// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     Oct 23 2022 18:16:08

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    led,
    usb_tx,
    trigger,
    rst_n,
    clk);

    output [7:0] led;
    output usb_tx;
    input trigger;
    input rst_n;
    input clk;

    wire N__3298;
    wire N__3297;
    wire N__3296;
    wire N__3287;
    wire N__3286;
    wire N__3285;
    wire N__3278;
    wire N__3277;
    wire N__3276;
    wire N__3269;
    wire N__3268;
    wire N__3267;
    wire N__3260;
    wire N__3259;
    wire N__3258;
    wire N__3251;
    wire N__3250;
    wire N__3249;
    wire N__3242;
    wire N__3241;
    wire N__3240;
    wire N__3233;
    wire N__3232;
    wire N__3231;
    wire N__3224;
    wire N__3223;
    wire N__3222;
    wire N__3215;
    wire N__3214;
    wire N__3213;
    wire N__3206;
    wire N__3205;
    wire N__3204;
    wire N__3197;
    wire N__3196;
    wire N__3195;
    wire N__3178;
    wire N__3175;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3160;
    wire N__3159;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3139;
    wire N__3138;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3128;
    wire N__3121;
    wire N__3120;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3097;
    wire N__3096;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3072;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3055;
    wire N__3052;
    wire N__3051;
    wire N__3048;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3024;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3007;
    wire N__3006;
    wire N__3003;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2986;
    wire N__2985;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2965;
    wire N__2962;
    wire N__2961;
    wire N__2958;
    wire N__2957;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2904;
    wire N__2903;
    wire N__2902;
    wire N__2901;
    wire N__2900;
    wire N__2899;
    wire N__2898;
    wire N__2897;
    wire N__2896;
    wire N__2895;
    wire N__2894;
    wire N__2893;
    wire N__2892;
    wire N__2891;
    wire N__2890;
    wire N__2889;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2819;
    wire N__2818;
    wire N__2815;
    wire N__2810;
    wire N__2807;
    wire N__2800;
    wire N__2797;
    wire N__2794;
    wire N__2791;
    wire N__2790;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2766;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2725;
    wire N__2724;
    wire N__2723;
    wire N__2720;
    wire N__2715;
    wire N__2714;
    wire N__2709;
    wire N__2706;
    wire N__2701;
    wire N__2698;
    wire N__2695;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2683;
    wire N__2682;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2665;
    wire N__2664;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2647;
    wire N__2646;
    wire N__2645;
    wire N__2642;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2626;
    wire N__2623;
    wire N__2622;
    wire N__2619;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2602;
    wire N__2601;
    wire N__2598;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2581;
    wire N__2580;
    wire N__2577;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2560;
    wire N__2559;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2539;
    wire N__2538;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2521;
    wire N__2520;
    wire N__2517;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2500;
    wire N__2499;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2482;
    wire N__2479;
    wire N__2476;
    wire N__2473;
    wire N__2470;
    wire N__2467;
    wire N__2464;
    wire N__2461;
    wire N__2460;
    wire N__2459;
    wire N__2452;
    wire N__2449;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2437;
    wire N__2436;
    wire N__2435;
    wire N__2434;
    wire N__2433;
    wire N__2430;
    wire N__2427;
    wire N__2426;
    wire N__2425;
    wire N__2424;
    wire N__2421;
    wire N__2420;
    wire N__2415;
    wire N__2412;
    wire N__2403;
    wire N__2398;
    wire N__2389;
    wire N__2388;
    wire N__2385;
    wire N__2384;
    wire N__2383;
    wire N__2382;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2376;
    wire N__2373;
    wire N__2366;
    wire N__2357;
    wire N__2350;
    wire N__2347;
    wire N__2344;
    wire N__2341;
    wire N__2338;
    wire N__2335;
    wire N__2332;
    wire N__2329;
    wire N__2328;
    wire N__2327;
    wire N__2324;
    wire N__2323;
    wire N__2318;
    wire N__2317;
    wire N__2316;
    wire N__2315;
    wire N__2314;
    wire N__2313;
    wire N__2312;
    wire N__2311;
    wire N__2310;
    wire N__2309;
    wire N__2306;
    wire N__2305;
    wire N__2304;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2287;
    wire N__2282;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire N__2266;
    wire N__2263;
    wire N__2242;
    wire N__2239;
    wire N__2238;
    wire N__2235;
    wire N__2234;
    wire N__2231;
    wire N__2230;
    wire N__2227;
    wire N__2224;
    wire N__2219;
    wire N__2212;
    wire N__2209;
    wire N__2206;
    wire N__2203;
    wire N__2200;
    wire N__2199;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2189;
    wire N__2184;
    wire N__2181;
    wire N__2176;
    wire N__2173;
    wire N__2170;
    wire N__2167;
    wire N__2164;
    wire N__2163;
    wire N__2162;
    wire N__2159;
    wire N__2156;
    wire N__2153;
    wire N__2146;
    wire N__2143;
    wire N__2140;
    wire N__2137;
    wire N__2134;
    wire N__2133;
    wire N__2130;
    wire N__2127;
    wire N__2122;
    wire N__2119;
    wire N__2116;
    wire N__2113;
    wire N__2110;
    wire N__2107;
    wire N__2104;
    wire N__2101;
    wire N__2098;
    wire N__2095;
    wire N__2092;
    wire N__2091;
    wire N__2090;
    wire N__2089;
    wire N__2088;
    wire N__2083;
    wire N__2080;
    wire N__2077;
    wire N__2074;
    wire N__2065;
    wire N__2064;
    wire N__2063;
    wire N__2062;
    wire N__2061;
    wire N__2058;
    wire N__2055;
    wire N__2050;
    wire N__2047;
    wire N__2044;
    wire N__2041;
    wire N__2032;
    wire N__2031;
    wire N__2030;
    wire N__2029;
    wire N__2026;
    wire N__2023;
    wire N__2020;
    wire N__2017;
    wire N__2008;
    wire N__2007;
    wire N__2006;
    wire N__2005;
    wire N__2004;
    wire N__2001;
    wire N__1998;
    wire N__1997;
    wire N__1994;
    wire N__1991;
    wire N__1988;
    wire N__1985;
    wire N__1982;
    wire N__1977;
    wire N__1966;
    wire N__1963;
    wire N__1960;
    wire N__1957;
    wire N__1954;
    wire N__1951;
    wire N__1948;
    wire N__1945;
    wire N__1942;
    wire N__1941;
    wire N__1938;
    wire N__1935;
    wire N__1932;
    wire N__1927;
    wire N__1924;
    wire N__1923;
    wire N__1922;
    wire N__1921;
    wire N__1920;
    wire N__1919;
    wire N__1918;
    wire N__1915;
    wire N__1908;
    wire N__1901;
    wire N__1894;
    wire N__1893;
    wire N__1890;
    wire N__1887;
    wire N__1882;
    wire N__1879;
    wire N__1876;
    wire N__1873;
    wire N__1872;
    wire N__1871;
    wire N__1870;
    wire N__1865;
    wire N__1860;
    wire N__1855;
    wire N__1852;
    wire N__1849;
    wire N__1848;
    wire N__1847;
    wire N__1846;
    wire N__1845;
    wire N__1842;
    wire N__1839;
    wire N__1834;
    wire N__1831;
    wire N__1822;
    wire N__1819;
    wire N__1816;
    wire N__1813;
    wire N__1810;
    wire N__1807;
    wire N__1804;
    wire N__1803;
    wire N__1802;
    wire N__1801;
    wire N__1800;
    wire N__1799;
    wire N__1796;
    wire N__1785;
    wire N__1780;
    wire N__1777;
    wire N__1774;
    wire N__1771;
    wire N__1768;
    wire N__1765;
    wire N__1764;
    wire N__1763;
    wire N__1762;
    wire N__1759;
    wire N__1752;
    wire N__1749;
    wire N__1746;
    wire N__1741;
    wire N__1738;
    wire N__1735;
    wire N__1732;
    wire N__1729;
    wire N__1726;
    wire N__1723;
    wire N__1722;
    wire N__1719;
    wire N__1716;
    wire N__1713;
    wire N__1708;
    wire N__1707;
    wire N__1704;
    wire N__1701;
    wire N__1696;
    wire N__1695;
    wire N__1692;
    wire N__1689;
    wire N__1686;
    wire N__1681;
    wire N__1678;
    wire N__1677;
    wire N__1674;
    wire N__1671;
    wire N__1666;
    wire N__1663;
    wire N__1660;
    wire N__1657;
    wire N__1656;
    wire N__1653;
    wire N__1650;
    wire N__1645;
    wire N__1642;
    wire N__1641;
    wire N__1638;
    wire N__1635;
    wire N__1630;
    wire N__1627;
    wire N__1626;
    wire N__1623;
    wire N__1620;
    wire N__1615;
    wire N__1612;
    wire N__1609;
    wire N__1606;
    wire N__1603;
    wire N__1600;
    wire N__1597;
    wire N__1594;
    wire N__1591;
    wire N__1588;
    wire N__1587;
    wire N__1586;
    wire N__1585;
    wire N__1582;
    wire N__1575;
    wire N__1572;
    wire N__1567;
    wire N__1564;
    wire N__1561;
    wire N__1558;
    wire N__1555;
    wire N__1552;
    wire N__1549;
    wire N__1546;
    wire N__1543;
    wire N__1540;
    wire N__1537;
    wire N__1536;
    wire N__1533;
    wire N__1530;
    wire N__1525;
    wire N__1524;
    wire N__1523;
    wire N__1522;
    wire N__1521;
    wire N__1516;
    wire N__1513;
    wire N__1510;
    wire N__1507;
    wire N__1498;
    wire N__1497;
    wire N__1496;
    wire N__1493;
    wire N__1490;
    wire N__1487;
    wire N__1484;
    wire N__1483;
    wire N__1480;
    wire N__1477;
    wire N__1474;
    wire N__1471;
    wire N__1470;
    wire N__1467;
    wire N__1460;
    wire N__1457;
    wire N__1450;
    wire N__1447;
    wire N__1444;
    wire N__1441;
    wire N__1438;
    wire N__1435;
    wire N__1432;
    wire N__1429;
    wire N__1426;
    wire N__1425;
    wire N__1424;
    wire N__1423;
    wire N__1414;
    wire N__1411;
    wire N__1408;
    wire N__1407;
    wire N__1404;
    wire N__1401;
    wire N__1396;
    wire N__1393;
    wire VCCG0;
    wire GNDG0;
    wire un1_M_count_q_ac0_1_cascade_;
    wire un1_M_count_q_ac0_1;
    wire click_dtct_out3_cascade_;
    wire un1_M_count_q_ac0_7_cascade_;
    wire click_dtct_out_d;
    wire click_dtct_out_d_cascade_;
    wire un1_M_count_q_ac0_7;
    wire \uart_tx.N_134_i_cascade_ ;
    wire \uart_tx.M_state_q_ns_0_o2_4_0_cascade_ ;
    wire \uart_tx.N_182_0_cascade_ ;
    wire \uart_tx.N_143_0_cascade_ ;
    wire uart_tx_N_185_cascade_;
    wire click_dtct_M_count_d6_0_1_cascade_;
    wire \uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_ ;
    wire uart_tx_N_187;
    wire un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_;
    wire un1_M_count_q_ac0_5_m2_0_a2_3;
    wire un1_M_count_q_ac0_5_m2_0_a2_3_cascade_;
    wire un1_M_count_q_ac0_out;
    wire click_dtct_out3;
    wire M_reset_cond_out_0;
    wire un1_M_count_q_axbxc7_1;
    wire \btn_cond.out_17_6_cascade_ ;
    wire \btn_cond.out_17_8 ;
    wire btn_cond_out_17_cascade_;
    wire click_dtct_out8;
    wire \btn_cond.out_17_7 ;
    wire \reset_cond.M_stage_qZ0Z_2 ;
    wire rst_n_c;
    wire \reset_cond.M_stage_qZ0Z_0 ;
    wire \reset_cond.M_stage_qZ0Z_1 ;
    wire \uart_tx.N_186_1_i ;
    wire \uart_tx.M_ctr_qZ0Z_0 ;
    wire bfn_15_22_0_;
    wire \uart_tx.M_ctr_qZ1Z_1 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_0 ;
    wire \uart_tx.M_ctr_qZ0Z_2 ;
    wire \uart_tx.M_ctr_q_RNO_0Z0Z_2 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_1 ;
    wire \uart_tx.M_ctr_qZ0Z_3 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_2 ;
    wire \uart_tx.M_ctr_qZ1Z_4 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_3 ;
    wire \uart_tx.M_ctr_qZ1Z_5 ;
    wire \uart_tx.M_ctr_q_RNO_0Z0Z_5 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_4 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_5 ;
    wire \uart_tx.N_134_i ;
    wire \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_ ;
    wire \uart_tx.N_182_0 ;
    wire \uart_tx.M_ctr_qZ0Z_6 ;
    wire \uart_tx.N_143_0 ;
    wire \uart_tx.M_bitCtr_qZ0Z_1 ;
    wire \uart_tx.M_txReg_q_RNOZ0Z_4_cascade_ ;
    wire \uart_tx.M_bitCtr_qZ1Z_0 ;
    wire \uart_tx.M_txReg_q_RNOZ0Z_2 ;
    wire \uart_tx.M_txReg_d_3_7_ns_1_cascade_ ;
    wire \uart_tx.M_txReg_q_RNOZ0Z_1 ;
    wire \uart_tx.M_bitCtr_qZ0Z_2 ;
    wire \uart_tx.M_txReg_q_RNOZ0Z_5 ;
    wire btn_cond_out_16_5;
    wire btn_cond_out_16_4;
    wire btn_cond_out_17;
    wire click_dtct_M_last_q;
    wire M_btn_cond_out_0_cascade_;
    wire bfn_15_25_0_;
    wire \btn_cond.un1_M_ctr_q_cry_0 ;
    wire \btn_cond.un1_M_ctr_q_cry_1 ;
    wire \btn_cond.un1_M_ctr_q_cry_2 ;
    wire \btn_cond.un1_M_ctr_q_cry_3 ;
    wire \btn_cond.un1_M_ctr_q_cry_4 ;
    wire \btn_cond.un1_M_ctr_q_cry_5 ;
    wire \btn_cond.un1_M_ctr_q_cry_6 ;
    wire \btn_cond.un1_M_ctr_q_cry_7 ;
    wire bfn_15_26_0_;
    wire \btn_cond.un1_M_ctr_q_cry_8 ;
    wire \btn_cond.un1_M_ctr_q_cry_9 ;
    wire \btn_cond.un1_M_ctr_q_cry_10 ;
    wire \btn_cond.un1_M_ctr_q_cry_11 ;
    wire \btn_cond.un1_M_ctr_q_cry_12 ;
    wire \btn_cond.un1_M_ctr_q_cry_13 ;
    wire \btn_cond.un1_M_ctr_q_cry_14 ;
    wire \btn_cond.un1_M_ctr_q_cry_15 ;
    wire bfn_15_27_0_;
    wire \btn_cond.un1_M_ctr_q_cry_16 ;
    wire \btn_cond.un1_M_ctr_q_cry_17 ;
    wire \btn_cond.un1_M_ctr_q_cry_18 ;
    wire \btn_cond.M_sync_out_i_g_0 ;
    wire \uart_tx.M_txReg_d_3 ;
    wire \uart_tx.M_state_qZ0Z_0 ;
    wire \uart_tx.M_state_qZ0Z_1 ;
    wire usb_tx_c;
    wire uart_tx_N_186_1;
    wire M_count_qZ0Z_0;
    wire \uart_tx.M_savedData_qZ0Z_0 ;
    wire M_count_qZ0Z_6;
    wire \uart_tx.M_savedData_qZ0Z_6 ;
    wire M_count_qZ0Z_4;
    wire \uart_tx.M_savedData_qZ0Z_4 ;
    wire M_count_qZ0Z_7;
    wire \uart_tx.M_savedData_qZ0Z_7 ;
    wire M_count_qZ0Z_2;
    wire \uart_tx.M_savedData_qZ0Z_2 ;
    wire M_count_qZ0Z_3;
    wire \uart_tx.M_savedData_qZ0Z_3 ;
    wire M_count_qZ0Z_1;
    wire \uart_tx.M_savedData_qZ0Z_1 ;
    wire M_count_qZ0Z_5;
    wire \uart_tx.M_savedData_qZ0Z_5 ;
    wire M_count_d6;
    wire \btn_cond.M_ctr_qZ0Z_6 ;
    wire \btn_cond.M_ctr_qZ0Z_5 ;
    wire \btn_cond.M_ctr_qZ0Z_4 ;
    wire \btn_cond.M_ctr_qZ0Z_7 ;
    wire \btn_cond.M_ctr_qZ0Z_11 ;
    wire \btn_cond.M_ctr_qZ0Z_8 ;
    wire \btn_cond.M_ctr_qZ0Z_10 ;
    wire \btn_cond.M_ctr_qZ0Z_9 ;
    wire \btn_cond.M_ctr_qZ0Z_15 ;
    wire \btn_cond.M_ctr_qZ0Z_14 ;
    wire \btn_cond.g0_13_cascade_ ;
    wire \btn_cond.g0_14 ;
    wire \btn_cond.g0_16_cascade_ ;
    wire \btn_cond.M_btn_cond_out_i_0 ;
    wire \btn_cond.M_ctr_qZ0Z_2 ;
    wire \btn_cond.M_ctr_qZ0Z_0 ;
    wire \btn_cond.M_ctr_qZ0Z_3 ;
    wire \btn_cond.M_ctr_qZ0Z_1 ;
    wire \btn_cond.g0_11 ;
    wire \btn_cond.M_ctr_qZ0Z_12 ;
    wire \btn_cond.M_ctr_qZ0Z_13 ;
    wire \btn_cond.g0_5 ;
    wire \btn_cond.M_ctr_qZ0Z_18 ;
    wire \btn_cond.M_ctr_qZ0Z_17 ;
    wire \btn_cond.M_ctr_qZ0Z_19 ;
    wire \btn_cond.M_ctr_qZ0Z_16 ;
    wire \btn_cond.g0_10 ;
    wire trigger_c;
    wire \btn_cond.sync.M_pipe_qZ0Z_0 ;
    wire clk_c_g;
    wire \btn_cond.sync.M_sync_out_0 ;
    wire \btn_cond.sync.M_sync_out_i_0 ;
    wire _gnd_net_;

    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3296),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__3298),
            .DIN(N__3297),
            .DOUT(N__3296),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__3298),
            .PADOUT(N__3297),
            .PADIN(N__3296),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__3287),
            .DIN(N__3286),
            .DOUT(N__3285),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__3287),
            .PADOUT(N__3286),
            .PADIN(N__3285),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__3278),
            .DIN(N__3277),
            .DOUT(N__3276),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__3278),
            .PADOUT(N__3277),
            .PADIN(N__3276),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__3269),
            .DIN(N__3268),
            .DOUT(N__3267),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__3269),
            .PADOUT(N__3268),
            .PADIN(N__3267),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__3260),
            .DIN(N__3259),
            .DOUT(N__3258),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__3260),
            .PADOUT(N__3259),
            .PADIN(N__3258),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__3251),
            .DIN(N__3250),
            .DOUT(N__3249),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__3251),
            .PADOUT(N__3250),
            .PADIN(N__3249),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__3242),
            .DIN(N__3241),
            .DOUT(N__3240),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__3242),
            .PADOUT(N__3241),
            .PADIN(N__3240),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__3233),
            .DIN(N__3232),
            .DOUT(N__3231),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__3233),
            .PADOUT(N__3232),
            .PADIN(N__3231),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__3224),
            .DIN(N__3223),
            .DOUT(N__3222),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__3224),
            .PADOUT(N__3223),
            .PADIN(N__3222),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__3215),
            .DIN(N__3214),
            .DOUT(N__3213),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__3215),
            .PADOUT(N__3214),
            .PADIN(N__3213),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD trigger_ibuf_iopad (
            .OE(N__3206),
            .DIN(N__3205),
            .DOUT(N__3204),
            .PACKAGEPIN(trigger));
    defparam trigger_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam trigger_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO trigger_ibuf_preio (
            .PADOEN(N__3206),
            .PADOUT(N__3205),
            .PADIN(N__3204),
            .CLOCKENABLE(),
            .DIN0(trigger_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD usb_tx_obuf_iopad (
            .OE(N__3197),
            .DIN(N__3196),
            .DOUT(N__3195),
            .PACKAGEPIN(usb_tx));
    defparam usb_tx_obuf_preio.NEG_TRIGGER=1'b0;
    defparam usb_tx_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO usb_tx_obuf_preio (
            .PADOEN(N__3197),
            .PADOUT(N__3196),
            .PADIN(N__3195),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2350),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__715 (
            .O(N__3178),
            .I(\btn_cond.g0_16_cascade_ ));
    CascadeMux I__714 (
            .O(N__3175),
            .I(N__3171));
    InMux I__713 (
            .O(N__3174),
            .I(N__3168));
    InMux I__712 (
            .O(N__3171),
            .I(N__3165));
    LocalMux I__711 (
            .O(N__3168),
            .I(\btn_cond.M_btn_cond_out_i_0 ));
    LocalMux I__710 (
            .O(N__3165),
            .I(\btn_cond.M_btn_cond_out_i_0 ));
    InMux I__709 (
            .O(N__3160),
            .I(N__3155));
    InMux I__708 (
            .O(N__3159),
            .I(N__3152));
    InMux I__707 (
            .O(N__3158),
            .I(N__3149));
    LocalMux I__706 (
            .O(N__3155),
            .I(N__3146));
    LocalMux I__705 (
            .O(N__3152),
            .I(\btn_cond.M_ctr_qZ0Z_2 ));
    LocalMux I__704 (
            .O(N__3149),
            .I(\btn_cond.M_ctr_qZ0Z_2 ));
    Odrv4 I__703 (
            .O(N__3146),
            .I(\btn_cond.M_ctr_qZ0Z_2 ));
    InMux I__702 (
            .O(N__3139),
            .I(N__3134));
    InMux I__701 (
            .O(N__3138),
            .I(N__3131));
    InMux I__700 (
            .O(N__3137),
            .I(N__3128));
    LocalMux I__699 (
            .O(N__3134),
            .I(\btn_cond.M_ctr_qZ0Z_0 ));
    LocalMux I__698 (
            .O(N__3131),
            .I(\btn_cond.M_ctr_qZ0Z_0 ));
    LocalMux I__697 (
            .O(N__3128),
            .I(\btn_cond.M_ctr_qZ0Z_0 ));
    CascadeMux I__696 (
            .O(N__3121),
            .I(N__3116));
    CascadeMux I__695 (
            .O(N__3120),
            .I(N__3113));
    InMux I__694 (
            .O(N__3119),
            .I(N__3110));
    InMux I__693 (
            .O(N__3116),
            .I(N__3107));
    InMux I__692 (
            .O(N__3113),
            .I(N__3104));
    LocalMux I__691 (
            .O(N__3110),
            .I(\btn_cond.M_ctr_qZ0Z_3 ));
    LocalMux I__690 (
            .O(N__3107),
            .I(\btn_cond.M_ctr_qZ0Z_3 ));
    LocalMux I__689 (
            .O(N__3104),
            .I(\btn_cond.M_ctr_qZ0Z_3 ));
    InMux I__688 (
            .O(N__3097),
            .I(N__3092));
    InMux I__687 (
            .O(N__3096),
            .I(N__3089));
    InMux I__686 (
            .O(N__3095),
            .I(N__3086));
    LocalMux I__685 (
            .O(N__3092),
            .I(\btn_cond.M_ctr_qZ0Z_1 ));
    LocalMux I__684 (
            .O(N__3089),
            .I(\btn_cond.M_ctr_qZ0Z_1 ));
    LocalMux I__683 (
            .O(N__3086),
            .I(\btn_cond.M_ctr_qZ0Z_1 ));
    InMux I__682 (
            .O(N__3079),
            .I(N__3076));
    LocalMux I__681 (
            .O(N__3076),
            .I(\btn_cond.g0_11 ));
    InMux I__680 (
            .O(N__3073),
            .I(N__3068));
    InMux I__679 (
            .O(N__3072),
            .I(N__3065));
    InMux I__678 (
            .O(N__3071),
            .I(N__3062));
    LocalMux I__677 (
            .O(N__3068),
            .I(\btn_cond.M_ctr_qZ0Z_12 ));
    LocalMux I__676 (
            .O(N__3065),
            .I(\btn_cond.M_ctr_qZ0Z_12 ));
    LocalMux I__675 (
            .O(N__3062),
            .I(\btn_cond.M_ctr_qZ0Z_12 ));
    InMux I__674 (
            .O(N__3055),
            .I(N__3052));
    LocalMux I__673 (
            .O(N__3052),
            .I(N__3048));
    InMux I__672 (
            .O(N__3051),
            .I(N__3044));
    Span4Mux_v I__671 (
            .O(N__3048),
            .I(N__3041));
    InMux I__670 (
            .O(N__3047),
            .I(N__3038));
    LocalMux I__669 (
            .O(N__3044),
            .I(\btn_cond.M_ctr_qZ0Z_13 ));
    Odrv4 I__668 (
            .O(N__3041),
            .I(\btn_cond.M_ctr_qZ0Z_13 ));
    LocalMux I__667 (
            .O(N__3038),
            .I(\btn_cond.M_ctr_qZ0Z_13 ));
    InMux I__666 (
            .O(N__3031),
            .I(N__3028));
    LocalMux I__665 (
            .O(N__3028),
            .I(\btn_cond.g0_5 ));
    InMux I__664 (
            .O(N__3025),
            .I(N__3020));
    InMux I__663 (
            .O(N__3024),
            .I(N__3017));
    InMux I__662 (
            .O(N__3023),
            .I(N__3014));
    LocalMux I__661 (
            .O(N__3020),
            .I(\btn_cond.M_ctr_qZ0Z_18 ));
    LocalMux I__660 (
            .O(N__3017),
            .I(\btn_cond.M_ctr_qZ0Z_18 ));
    LocalMux I__659 (
            .O(N__3014),
            .I(\btn_cond.M_ctr_qZ0Z_18 ));
    InMux I__658 (
            .O(N__3007),
            .I(N__3003));
    InMux I__657 (
            .O(N__3006),
            .I(N__2999));
    LocalMux I__656 (
            .O(N__3003),
            .I(N__2996));
    InMux I__655 (
            .O(N__3002),
            .I(N__2993));
    LocalMux I__654 (
            .O(N__2999),
            .I(\btn_cond.M_ctr_qZ0Z_17 ));
    Odrv4 I__653 (
            .O(N__2996),
            .I(\btn_cond.M_ctr_qZ0Z_17 ));
    LocalMux I__652 (
            .O(N__2993),
            .I(\btn_cond.M_ctr_qZ0Z_17 ));
    CascadeMux I__651 (
            .O(N__2986),
            .I(N__2981));
    InMux I__650 (
            .O(N__2985),
            .I(N__2978));
    InMux I__649 (
            .O(N__2984),
            .I(N__2975));
    InMux I__648 (
            .O(N__2981),
            .I(N__2972));
    LocalMux I__647 (
            .O(N__2978),
            .I(\btn_cond.M_ctr_qZ0Z_19 ));
    LocalMux I__646 (
            .O(N__2975),
            .I(\btn_cond.M_ctr_qZ0Z_19 ));
    LocalMux I__645 (
            .O(N__2972),
            .I(\btn_cond.M_ctr_qZ0Z_19 ));
    CascadeMux I__644 (
            .O(N__2965),
            .I(N__2962));
    InMux I__643 (
            .O(N__2962),
            .I(N__2958));
    InMux I__642 (
            .O(N__2961),
            .I(N__2954));
    LocalMux I__641 (
            .O(N__2958),
            .I(N__2951));
    InMux I__640 (
            .O(N__2957),
            .I(N__2948));
    LocalMux I__639 (
            .O(N__2954),
            .I(\btn_cond.M_ctr_qZ0Z_16 ));
    Odrv4 I__638 (
            .O(N__2951),
            .I(\btn_cond.M_ctr_qZ0Z_16 ));
    LocalMux I__637 (
            .O(N__2948),
            .I(\btn_cond.M_ctr_qZ0Z_16 ));
    InMux I__636 (
            .O(N__2941),
            .I(N__2938));
    LocalMux I__635 (
            .O(N__2938),
            .I(\btn_cond.g0_10 ));
    InMux I__634 (
            .O(N__2935),
            .I(N__2932));
    LocalMux I__633 (
            .O(N__2932),
            .I(N__2929));
    Span4Mux_v I__632 (
            .O(N__2929),
            .I(N__2926));
    Sp12to4 I__631 (
            .O(N__2926),
            .I(N__2923));
    Span12Mux_h I__630 (
            .O(N__2923),
            .I(N__2920));
    Span12Mux_v I__629 (
            .O(N__2920),
            .I(N__2917));
    Span12Mux_v I__628 (
            .O(N__2917),
            .I(N__2914));
    Odrv12 I__627 (
            .O(N__2914),
            .I(trigger_c));
    InMux I__626 (
            .O(N__2911),
            .I(N__2908));
    LocalMux I__625 (
            .O(N__2908),
            .I(\btn_cond.sync.M_pipe_qZ0Z_0 ));
    ClkMux I__624 (
            .O(N__2905),
            .I(N__2854));
    ClkMux I__623 (
            .O(N__2904),
            .I(N__2854));
    ClkMux I__622 (
            .O(N__2903),
            .I(N__2854));
    ClkMux I__621 (
            .O(N__2902),
            .I(N__2854));
    ClkMux I__620 (
            .O(N__2901),
            .I(N__2854));
    ClkMux I__619 (
            .O(N__2900),
            .I(N__2854));
    ClkMux I__618 (
            .O(N__2899),
            .I(N__2854));
    ClkMux I__617 (
            .O(N__2898),
            .I(N__2854));
    ClkMux I__616 (
            .O(N__2897),
            .I(N__2854));
    ClkMux I__615 (
            .O(N__2896),
            .I(N__2854));
    ClkMux I__614 (
            .O(N__2895),
            .I(N__2854));
    ClkMux I__613 (
            .O(N__2894),
            .I(N__2854));
    ClkMux I__612 (
            .O(N__2893),
            .I(N__2854));
    ClkMux I__611 (
            .O(N__2892),
            .I(N__2854));
    ClkMux I__610 (
            .O(N__2891),
            .I(N__2854));
    ClkMux I__609 (
            .O(N__2890),
            .I(N__2854));
    ClkMux I__608 (
            .O(N__2889),
            .I(N__2854));
    GlobalMux I__607 (
            .O(N__2854),
            .I(N__2851));
    gio2CtrlBuf I__606 (
            .O(N__2851),
            .I(clk_c_g));
    InMux I__605 (
            .O(N__2848),
            .I(N__2845));
    LocalMux I__604 (
            .O(N__2845),
            .I(\btn_cond.sync.M_sync_out_0 ));
    IoInMux I__603 (
            .O(N__2842),
            .I(N__2839));
    LocalMux I__602 (
            .O(N__2839),
            .I(\btn_cond.sync.M_sync_out_i_0 ));
    InMux I__601 (
            .O(N__2836),
            .I(N__2833));
    LocalMux I__600 (
            .O(N__2833),
            .I(N__2830));
    Odrv4 I__599 (
            .O(N__2830),
            .I(\uart_tx.M_savedData_qZ0Z_7 ));
    InMux I__598 (
            .O(N__2827),
            .I(N__2823));
    CascadeMux I__597 (
            .O(N__2826),
            .I(N__2820));
    LocalMux I__596 (
            .O(N__2823),
            .I(N__2815));
    InMux I__595 (
            .O(N__2820),
            .I(N__2810));
    InMux I__594 (
            .O(N__2819),
            .I(N__2810));
    InMux I__593 (
            .O(N__2818),
            .I(N__2807));
    Odrv4 I__592 (
            .O(N__2815),
            .I(M_count_qZ0Z_2));
    LocalMux I__591 (
            .O(N__2810),
            .I(M_count_qZ0Z_2));
    LocalMux I__590 (
            .O(N__2807),
            .I(M_count_qZ0Z_2));
    InMux I__589 (
            .O(N__2800),
            .I(N__2797));
    LocalMux I__588 (
            .O(N__2797),
            .I(\uart_tx.M_savedData_qZ0Z_2 ));
    InMux I__587 (
            .O(N__2794),
            .I(N__2791));
    LocalMux I__586 (
            .O(N__2791),
            .I(N__2786));
    InMux I__585 (
            .O(N__2790),
            .I(N__2783));
    InMux I__584 (
            .O(N__2789),
            .I(N__2780));
    Odrv4 I__583 (
            .O(N__2786),
            .I(M_count_qZ0Z_3));
    LocalMux I__582 (
            .O(N__2783),
            .I(M_count_qZ0Z_3));
    LocalMux I__581 (
            .O(N__2780),
            .I(M_count_qZ0Z_3));
    InMux I__580 (
            .O(N__2773),
            .I(N__2770));
    LocalMux I__579 (
            .O(N__2770),
            .I(\uart_tx.M_savedData_qZ0Z_3 ));
    InMux I__578 (
            .O(N__2767),
            .I(N__2762));
    CascadeMux I__577 (
            .O(N__2766),
            .I(N__2759));
    InMux I__576 (
            .O(N__2765),
            .I(N__2756));
    LocalMux I__575 (
            .O(N__2762),
            .I(N__2752));
    InMux I__574 (
            .O(N__2759),
            .I(N__2749));
    LocalMux I__573 (
            .O(N__2756),
            .I(N__2746));
    InMux I__572 (
            .O(N__2755),
            .I(N__2743));
    Odrv4 I__571 (
            .O(N__2752),
            .I(M_count_qZ0Z_1));
    LocalMux I__570 (
            .O(N__2749),
            .I(M_count_qZ0Z_1));
    Odrv4 I__569 (
            .O(N__2746),
            .I(M_count_qZ0Z_1));
    LocalMux I__568 (
            .O(N__2743),
            .I(M_count_qZ0Z_1));
    InMux I__567 (
            .O(N__2734),
            .I(N__2731));
    LocalMux I__566 (
            .O(N__2731),
            .I(\uart_tx.M_savedData_qZ0Z_1 ));
    InMux I__565 (
            .O(N__2728),
            .I(N__2725));
    LocalMux I__564 (
            .O(N__2725),
            .I(N__2720));
    InMux I__563 (
            .O(N__2724),
            .I(N__2715));
    InMux I__562 (
            .O(N__2723),
            .I(N__2715));
    Span4Mux_h I__561 (
            .O(N__2720),
            .I(N__2709));
    LocalMux I__560 (
            .O(N__2715),
            .I(N__2709));
    InMux I__559 (
            .O(N__2714),
            .I(N__2706));
    Odrv4 I__558 (
            .O(N__2709),
            .I(M_count_qZ0Z_5));
    LocalMux I__557 (
            .O(N__2706),
            .I(M_count_qZ0Z_5));
    InMux I__556 (
            .O(N__2701),
            .I(N__2698));
    LocalMux I__555 (
            .O(N__2698),
            .I(\uart_tx.M_savedData_qZ0Z_5 ));
    CEMux I__554 (
            .O(N__2695),
            .I(N__2691));
    CEMux I__553 (
            .O(N__2694),
            .I(N__2688));
    LocalMux I__552 (
            .O(N__2691),
            .I(M_count_d6));
    LocalMux I__551 (
            .O(N__2688),
            .I(M_count_d6));
    InMux I__550 (
            .O(N__2683),
            .I(N__2678));
    InMux I__549 (
            .O(N__2682),
            .I(N__2675));
    InMux I__548 (
            .O(N__2681),
            .I(N__2672));
    LocalMux I__547 (
            .O(N__2678),
            .I(\btn_cond.M_ctr_qZ0Z_6 ));
    LocalMux I__546 (
            .O(N__2675),
            .I(\btn_cond.M_ctr_qZ0Z_6 ));
    LocalMux I__545 (
            .O(N__2672),
            .I(\btn_cond.M_ctr_qZ0Z_6 ));
    InMux I__544 (
            .O(N__2665),
            .I(N__2660));
    InMux I__543 (
            .O(N__2664),
            .I(N__2657));
    InMux I__542 (
            .O(N__2663),
            .I(N__2654));
    LocalMux I__541 (
            .O(N__2660),
            .I(\btn_cond.M_ctr_qZ0Z_5 ));
    LocalMux I__540 (
            .O(N__2657),
            .I(\btn_cond.M_ctr_qZ0Z_5 ));
    LocalMux I__539 (
            .O(N__2654),
            .I(\btn_cond.M_ctr_qZ0Z_5 ));
    CascadeMux I__538 (
            .O(N__2647),
            .I(N__2642));
    InMux I__537 (
            .O(N__2646),
            .I(N__2639));
    InMux I__536 (
            .O(N__2645),
            .I(N__2636));
    InMux I__535 (
            .O(N__2642),
            .I(N__2633));
    LocalMux I__534 (
            .O(N__2639),
            .I(\btn_cond.M_ctr_qZ0Z_4 ));
    LocalMux I__533 (
            .O(N__2636),
            .I(\btn_cond.M_ctr_qZ0Z_4 ));
    LocalMux I__532 (
            .O(N__2633),
            .I(\btn_cond.M_ctr_qZ0Z_4 ));
    CascadeMux I__531 (
            .O(N__2626),
            .I(N__2623));
    InMux I__530 (
            .O(N__2623),
            .I(N__2619));
    InMux I__529 (
            .O(N__2622),
            .I(N__2615));
    LocalMux I__528 (
            .O(N__2619),
            .I(N__2612));
    InMux I__527 (
            .O(N__2618),
            .I(N__2609));
    LocalMux I__526 (
            .O(N__2615),
            .I(\btn_cond.M_ctr_qZ0Z_7 ));
    Odrv12 I__525 (
            .O(N__2612),
            .I(\btn_cond.M_ctr_qZ0Z_7 ));
    LocalMux I__524 (
            .O(N__2609),
            .I(\btn_cond.M_ctr_qZ0Z_7 ));
    InMux I__523 (
            .O(N__2602),
            .I(N__2598));
    InMux I__522 (
            .O(N__2601),
            .I(N__2594));
    LocalMux I__521 (
            .O(N__2598),
            .I(N__2591));
    InMux I__520 (
            .O(N__2597),
            .I(N__2588));
    LocalMux I__519 (
            .O(N__2594),
            .I(\btn_cond.M_ctr_qZ0Z_11 ));
    Odrv4 I__518 (
            .O(N__2591),
            .I(\btn_cond.M_ctr_qZ0Z_11 ));
    LocalMux I__517 (
            .O(N__2588),
            .I(\btn_cond.M_ctr_qZ0Z_11 ));
    CascadeMux I__516 (
            .O(N__2581),
            .I(N__2577));
    InMux I__515 (
            .O(N__2580),
            .I(N__2573));
    InMux I__514 (
            .O(N__2577),
            .I(N__2570));
    InMux I__513 (
            .O(N__2576),
            .I(N__2567));
    LocalMux I__512 (
            .O(N__2573),
            .I(\btn_cond.M_ctr_qZ0Z_8 ));
    LocalMux I__511 (
            .O(N__2570),
            .I(\btn_cond.M_ctr_qZ0Z_8 ));
    LocalMux I__510 (
            .O(N__2567),
            .I(\btn_cond.M_ctr_qZ0Z_8 ));
    CascadeMux I__509 (
            .O(N__2560),
            .I(N__2555));
    InMux I__508 (
            .O(N__2559),
            .I(N__2552));
    InMux I__507 (
            .O(N__2558),
            .I(N__2549));
    InMux I__506 (
            .O(N__2555),
            .I(N__2546));
    LocalMux I__505 (
            .O(N__2552),
            .I(\btn_cond.M_ctr_qZ0Z_10 ));
    LocalMux I__504 (
            .O(N__2549),
            .I(\btn_cond.M_ctr_qZ0Z_10 ));
    LocalMux I__503 (
            .O(N__2546),
            .I(\btn_cond.M_ctr_qZ0Z_10 ));
    InMux I__502 (
            .O(N__2539),
            .I(N__2534));
    InMux I__501 (
            .O(N__2538),
            .I(N__2531));
    InMux I__500 (
            .O(N__2537),
            .I(N__2528));
    LocalMux I__499 (
            .O(N__2534),
            .I(\btn_cond.M_ctr_qZ0Z_9 ));
    LocalMux I__498 (
            .O(N__2531),
            .I(\btn_cond.M_ctr_qZ0Z_9 ));
    LocalMux I__497 (
            .O(N__2528),
            .I(\btn_cond.M_ctr_qZ0Z_9 ));
    CascadeMux I__496 (
            .O(N__2521),
            .I(N__2517));
    InMux I__495 (
            .O(N__2520),
            .I(N__2513));
    InMux I__494 (
            .O(N__2517),
            .I(N__2510));
    InMux I__493 (
            .O(N__2516),
            .I(N__2507));
    LocalMux I__492 (
            .O(N__2513),
            .I(\btn_cond.M_ctr_qZ0Z_15 ));
    LocalMux I__491 (
            .O(N__2510),
            .I(\btn_cond.M_ctr_qZ0Z_15 ));
    LocalMux I__490 (
            .O(N__2507),
            .I(\btn_cond.M_ctr_qZ0Z_15 ));
    InMux I__489 (
            .O(N__2500),
            .I(N__2495));
    InMux I__488 (
            .O(N__2499),
            .I(N__2492));
    InMux I__487 (
            .O(N__2498),
            .I(N__2489));
    LocalMux I__486 (
            .O(N__2495),
            .I(\btn_cond.M_ctr_qZ0Z_14 ));
    LocalMux I__485 (
            .O(N__2492),
            .I(\btn_cond.M_ctr_qZ0Z_14 ));
    LocalMux I__484 (
            .O(N__2489),
            .I(\btn_cond.M_ctr_qZ0Z_14 ));
    CascadeMux I__483 (
            .O(N__2482),
            .I(\btn_cond.g0_13_cascade_ ));
    InMux I__482 (
            .O(N__2479),
            .I(N__2476));
    LocalMux I__481 (
            .O(N__2476),
            .I(\btn_cond.g0_14 ));
    InMux I__480 (
            .O(N__2473),
            .I(bfn_15_27_0_));
    InMux I__479 (
            .O(N__2470),
            .I(\btn_cond.un1_M_ctr_q_cry_16 ));
    InMux I__478 (
            .O(N__2467),
            .I(\btn_cond.un1_M_ctr_q_cry_17 ));
    InMux I__477 (
            .O(N__2464),
            .I(\btn_cond.un1_M_ctr_q_cry_18 ));
    SRMux I__476 (
            .O(N__2461),
            .I(N__2452));
    SRMux I__475 (
            .O(N__2460),
            .I(N__2452));
    SRMux I__474 (
            .O(N__2459),
            .I(N__2452));
    GlobalMux I__473 (
            .O(N__2452),
            .I(N__2449));
    gio2CtrlBuf I__472 (
            .O(N__2449),
            .I(\btn_cond.M_sync_out_i_g_0 ));
    InMux I__471 (
            .O(N__2446),
            .I(N__2443));
    LocalMux I__470 (
            .O(N__2443),
            .I(\uart_tx.M_txReg_d_3 ));
    InMux I__469 (
            .O(N__2440),
            .I(N__2437));
    LocalMux I__468 (
            .O(N__2437),
            .I(N__2430));
    CascadeMux I__467 (
            .O(N__2436),
            .I(N__2427));
    CascadeMux I__466 (
            .O(N__2435),
            .I(N__2421));
    InMux I__465 (
            .O(N__2434),
            .I(N__2415));
    InMux I__464 (
            .O(N__2433),
            .I(N__2415));
    Span4Mux_h I__463 (
            .O(N__2430),
            .I(N__2412));
    InMux I__462 (
            .O(N__2427),
            .I(N__2403));
    InMux I__461 (
            .O(N__2426),
            .I(N__2403));
    InMux I__460 (
            .O(N__2425),
            .I(N__2403));
    InMux I__459 (
            .O(N__2424),
            .I(N__2403));
    InMux I__458 (
            .O(N__2421),
            .I(N__2398));
    InMux I__457 (
            .O(N__2420),
            .I(N__2398));
    LocalMux I__456 (
            .O(N__2415),
            .I(\uart_tx.M_state_qZ0Z_0 ));
    Odrv4 I__455 (
            .O(N__2412),
            .I(\uart_tx.M_state_qZ0Z_0 ));
    LocalMux I__454 (
            .O(N__2403),
            .I(\uart_tx.M_state_qZ0Z_0 ));
    LocalMux I__453 (
            .O(N__2398),
            .I(\uart_tx.M_state_qZ0Z_0 ));
    InMux I__452 (
            .O(N__2389),
            .I(N__2385));
    CascadeMux I__451 (
            .O(N__2388),
            .I(N__2379));
    LocalMux I__450 (
            .O(N__2385),
            .I(N__2373));
    InMux I__449 (
            .O(N__2384),
            .I(N__2366));
    InMux I__448 (
            .O(N__2383),
            .I(N__2366));
    InMux I__447 (
            .O(N__2382),
            .I(N__2366));
    InMux I__446 (
            .O(N__2379),
            .I(N__2357));
    InMux I__445 (
            .O(N__2378),
            .I(N__2357));
    InMux I__444 (
            .O(N__2377),
            .I(N__2357));
    InMux I__443 (
            .O(N__2376),
            .I(N__2357));
    Odrv4 I__442 (
            .O(N__2373),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    LocalMux I__441 (
            .O(N__2366),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    LocalMux I__440 (
            .O(N__2357),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    IoInMux I__439 (
            .O(N__2350),
            .I(N__2347));
    LocalMux I__438 (
            .O(N__2347),
            .I(N__2344));
    Span4Mux_s0_v I__437 (
            .O(N__2344),
            .I(N__2341));
    Sp12to4 I__436 (
            .O(N__2341),
            .I(N__2338));
    Span12Mux_h I__435 (
            .O(N__2338),
            .I(N__2335));
    Span12Mux_v I__434 (
            .O(N__2335),
            .I(N__2332));
    Odrv12 I__433 (
            .O(N__2332),
            .I(usb_tx_c));
    SRMux I__432 (
            .O(N__2329),
            .I(N__2324));
    InMux I__431 (
            .O(N__2328),
            .I(N__2318));
    InMux I__430 (
            .O(N__2327),
            .I(N__2318));
    LocalMux I__429 (
            .O(N__2324),
            .I(N__2306));
    InMux I__428 (
            .O(N__2323),
            .I(N__2300));
    LocalMux I__427 (
            .O(N__2318),
            .I(N__2297));
    InMux I__426 (
            .O(N__2317),
            .I(N__2294));
    InMux I__425 (
            .O(N__2316),
            .I(N__2287));
    InMux I__424 (
            .O(N__2315),
            .I(N__2287));
    InMux I__423 (
            .O(N__2314),
            .I(N__2287));
    InMux I__422 (
            .O(N__2313),
            .I(N__2282));
    InMux I__421 (
            .O(N__2312),
            .I(N__2282));
    InMux I__420 (
            .O(N__2311),
            .I(N__2275));
    InMux I__419 (
            .O(N__2310),
            .I(N__2275));
    InMux I__418 (
            .O(N__2309),
            .I(N__2275));
    Span4Mux_h I__417 (
            .O(N__2306),
            .I(N__2272));
    InMux I__416 (
            .O(N__2305),
            .I(N__2269));
    InMux I__415 (
            .O(N__2304),
            .I(N__2266));
    InMux I__414 (
            .O(N__2303),
            .I(N__2263));
    LocalMux I__413 (
            .O(N__2300),
            .I(uart_tx_N_186_1));
    Odrv4 I__412 (
            .O(N__2297),
            .I(uart_tx_N_186_1));
    LocalMux I__411 (
            .O(N__2294),
            .I(uart_tx_N_186_1));
    LocalMux I__410 (
            .O(N__2287),
            .I(uart_tx_N_186_1));
    LocalMux I__409 (
            .O(N__2282),
            .I(uart_tx_N_186_1));
    LocalMux I__408 (
            .O(N__2275),
            .I(uart_tx_N_186_1));
    Odrv4 I__407 (
            .O(N__2272),
            .I(uart_tx_N_186_1));
    LocalMux I__406 (
            .O(N__2269),
            .I(uart_tx_N_186_1));
    LocalMux I__405 (
            .O(N__2266),
            .I(uart_tx_N_186_1));
    LocalMux I__404 (
            .O(N__2263),
            .I(uart_tx_N_186_1));
    InMux I__403 (
            .O(N__2242),
            .I(N__2239));
    LocalMux I__402 (
            .O(N__2239),
            .I(N__2235));
    CascadeMux I__401 (
            .O(N__2238),
            .I(N__2231));
    Span4Mux_v I__400 (
            .O(N__2235),
            .I(N__2227));
    InMux I__399 (
            .O(N__2234),
            .I(N__2224));
    InMux I__398 (
            .O(N__2231),
            .I(N__2219));
    InMux I__397 (
            .O(N__2230),
            .I(N__2219));
    Odrv4 I__396 (
            .O(N__2227),
            .I(M_count_qZ0Z_0));
    LocalMux I__395 (
            .O(N__2224),
            .I(M_count_qZ0Z_0));
    LocalMux I__394 (
            .O(N__2219),
            .I(M_count_qZ0Z_0));
    InMux I__393 (
            .O(N__2212),
            .I(N__2209));
    LocalMux I__392 (
            .O(N__2209),
            .I(N__2206));
    Odrv4 I__391 (
            .O(N__2206),
            .I(\uart_tx.M_savedData_qZ0Z_0 ));
    InMux I__390 (
            .O(N__2203),
            .I(N__2200));
    LocalMux I__389 (
            .O(N__2200),
            .I(N__2195));
    InMux I__388 (
            .O(N__2199),
            .I(N__2192));
    InMux I__387 (
            .O(N__2198),
            .I(N__2189));
    Span4Mux_v I__386 (
            .O(N__2195),
            .I(N__2184));
    LocalMux I__385 (
            .O(N__2192),
            .I(N__2184));
    LocalMux I__384 (
            .O(N__2189),
            .I(N__2181));
    Odrv4 I__383 (
            .O(N__2184),
            .I(M_count_qZ0Z_6));
    Odrv4 I__382 (
            .O(N__2181),
            .I(M_count_qZ0Z_6));
    InMux I__381 (
            .O(N__2176),
            .I(N__2173));
    LocalMux I__380 (
            .O(N__2173),
            .I(\uart_tx.M_savedData_qZ0Z_6 ));
    InMux I__379 (
            .O(N__2170),
            .I(N__2167));
    LocalMux I__378 (
            .O(N__2167),
            .I(N__2164));
    Span4Mux_h I__377 (
            .O(N__2164),
            .I(N__2159));
    InMux I__376 (
            .O(N__2163),
            .I(N__2156));
    InMux I__375 (
            .O(N__2162),
            .I(N__2153));
    Odrv4 I__374 (
            .O(N__2159),
            .I(M_count_qZ0Z_4));
    LocalMux I__373 (
            .O(N__2156),
            .I(M_count_qZ0Z_4));
    LocalMux I__372 (
            .O(N__2153),
            .I(M_count_qZ0Z_4));
    InMux I__371 (
            .O(N__2146),
            .I(N__2143));
    LocalMux I__370 (
            .O(N__2143),
            .I(\uart_tx.M_savedData_qZ0Z_4 ));
    InMux I__369 (
            .O(N__2140),
            .I(N__2137));
    LocalMux I__368 (
            .O(N__2137),
            .I(N__2134));
    Span4Mux_v I__367 (
            .O(N__2134),
            .I(N__2130));
    InMux I__366 (
            .O(N__2133),
            .I(N__2127));
    Odrv4 I__365 (
            .O(N__2130),
            .I(M_count_qZ0Z_7));
    LocalMux I__364 (
            .O(N__2127),
            .I(M_count_qZ0Z_7));
    InMux I__363 (
            .O(N__2122),
            .I(\btn_cond.un1_M_ctr_q_cry_6 ));
    InMux I__362 (
            .O(N__2119),
            .I(bfn_15_26_0_));
    InMux I__361 (
            .O(N__2116),
            .I(\btn_cond.un1_M_ctr_q_cry_8 ));
    InMux I__360 (
            .O(N__2113),
            .I(\btn_cond.un1_M_ctr_q_cry_9 ));
    InMux I__359 (
            .O(N__2110),
            .I(\btn_cond.un1_M_ctr_q_cry_10 ));
    InMux I__358 (
            .O(N__2107),
            .I(\btn_cond.un1_M_ctr_q_cry_11 ));
    InMux I__357 (
            .O(N__2104),
            .I(\btn_cond.un1_M_ctr_q_cry_12 ));
    InMux I__356 (
            .O(N__2101),
            .I(\btn_cond.un1_M_ctr_q_cry_13 ));
    InMux I__355 (
            .O(N__2098),
            .I(\btn_cond.un1_M_ctr_q_cry_14 ));
    CascadeMux I__354 (
            .O(N__2095),
            .I(N__2092));
    InMux I__353 (
            .O(N__2092),
            .I(N__2083));
    InMux I__352 (
            .O(N__2091),
            .I(N__2083));
    InMux I__351 (
            .O(N__2090),
            .I(N__2080));
    InMux I__350 (
            .O(N__2089),
            .I(N__2077));
    InMux I__349 (
            .O(N__2088),
            .I(N__2074));
    LocalMux I__348 (
            .O(N__2083),
            .I(btn_cond_out_16_5));
    LocalMux I__347 (
            .O(N__2080),
            .I(btn_cond_out_16_5));
    LocalMux I__346 (
            .O(N__2077),
            .I(btn_cond_out_16_5));
    LocalMux I__345 (
            .O(N__2074),
            .I(btn_cond_out_16_5));
    InMux I__344 (
            .O(N__2065),
            .I(N__2058));
    InMux I__343 (
            .O(N__2064),
            .I(N__2055));
    InMux I__342 (
            .O(N__2063),
            .I(N__2050));
    InMux I__341 (
            .O(N__2062),
            .I(N__2050));
    InMux I__340 (
            .O(N__2061),
            .I(N__2047));
    LocalMux I__339 (
            .O(N__2058),
            .I(N__2044));
    LocalMux I__338 (
            .O(N__2055),
            .I(N__2041));
    LocalMux I__337 (
            .O(N__2050),
            .I(btn_cond_out_16_4));
    LocalMux I__336 (
            .O(N__2047),
            .I(btn_cond_out_16_4));
    Odrv4 I__335 (
            .O(N__2044),
            .I(btn_cond_out_16_4));
    Odrv4 I__334 (
            .O(N__2041),
            .I(btn_cond_out_16_4));
    InMux I__333 (
            .O(N__2032),
            .I(N__2026));
    InMux I__332 (
            .O(N__2031),
            .I(N__2023));
    InMux I__331 (
            .O(N__2030),
            .I(N__2020));
    InMux I__330 (
            .O(N__2029),
            .I(N__2017));
    LocalMux I__329 (
            .O(N__2026),
            .I(btn_cond_out_17));
    LocalMux I__328 (
            .O(N__2023),
            .I(btn_cond_out_17));
    LocalMux I__327 (
            .O(N__2020),
            .I(btn_cond_out_17));
    LocalMux I__326 (
            .O(N__2017),
            .I(btn_cond_out_17));
    CascadeMux I__325 (
            .O(N__2008),
            .I(N__2001));
    CascadeMux I__324 (
            .O(N__2007),
            .I(N__1998));
    CascadeMux I__323 (
            .O(N__2006),
            .I(N__1994));
    InMux I__322 (
            .O(N__2005),
            .I(N__1991));
    InMux I__321 (
            .O(N__2004),
            .I(N__1988));
    InMux I__320 (
            .O(N__2001),
            .I(N__1985));
    InMux I__319 (
            .O(N__1998),
            .I(N__1982));
    InMux I__318 (
            .O(N__1997),
            .I(N__1977));
    InMux I__317 (
            .O(N__1994),
            .I(N__1977));
    LocalMux I__316 (
            .O(N__1991),
            .I(click_dtct_M_last_q));
    LocalMux I__315 (
            .O(N__1988),
            .I(click_dtct_M_last_q));
    LocalMux I__314 (
            .O(N__1985),
            .I(click_dtct_M_last_q));
    LocalMux I__313 (
            .O(N__1982),
            .I(click_dtct_M_last_q));
    LocalMux I__312 (
            .O(N__1977),
            .I(click_dtct_M_last_q));
    CascadeMux I__311 (
            .O(N__1966),
            .I(M_btn_cond_out_0_cascade_));
    InMux I__310 (
            .O(N__1963),
            .I(\btn_cond.un1_M_ctr_q_cry_0 ));
    InMux I__309 (
            .O(N__1960),
            .I(\btn_cond.un1_M_ctr_q_cry_1 ));
    InMux I__308 (
            .O(N__1957),
            .I(\btn_cond.un1_M_ctr_q_cry_2 ));
    InMux I__307 (
            .O(N__1954),
            .I(\btn_cond.un1_M_ctr_q_cry_3 ));
    InMux I__306 (
            .O(N__1951),
            .I(\btn_cond.un1_M_ctr_q_cry_4 ));
    InMux I__305 (
            .O(N__1948),
            .I(\btn_cond.un1_M_ctr_q_cry_5 ));
    InMux I__304 (
            .O(N__1945),
            .I(\uart_tx.un1_M_ctr_q_3_cry_5 ));
    CascadeMux I__303 (
            .O(N__1942),
            .I(N__1938));
    InMux I__302 (
            .O(N__1941),
            .I(N__1935));
    InMux I__301 (
            .O(N__1938),
            .I(N__1932));
    LocalMux I__300 (
            .O(N__1935),
            .I(\uart_tx.N_134_i ));
    LocalMux I__299 (
            .O(N__1932),
            .I(\uart_tx.N_134_i ));
    CascadeMux I__298 (
            .O(N__1927),
            .I(\uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_ ));
    InMux I__297 (
            .O(N__1924),
            .I(N__1915));
    InMux I__296 (
            .O(N__1923),
            .I(N__1908));
    InMux I__295 (
            .O(N__1922),
            .I(N__1908));
    InMux I__294 (
            .O(N__1921),
            .I(N__1908));
    InMux I__293 (
            .O(N__1920),
            .I(N__1901));
    InMux I__292 (
            .O(N__1919),
            .I(N__1901));
    InMux I__291 (
            .O(N__1918),
            .I(N__1901));
    LocalMux I__290 (
            .O(N__1915),
            .I(\uart_tx.N_182_0 ));
    LocalMux I__289 (
            .O(N__1908),
            .I(\uart_tx.N_182_0 ));
    LocalMux I__288 (
            .O(N__1901),
            .I(\uart_tx.N_182_0 ));
    InMux I__287 (
            .O(N__1894),
            .I(N__1890));
    InMux I__286 (
            .O(N__1893),
            .I(N__1887));
    LocalMux I__285 (
            .O(N__1890),
            .I(\uart_tx.M_ctr_qZ0Z_6 ));
    LocalMux I__284 (
            .O(N__1887),
            .I(\uart_tx.M_ctr_qZ0Z_6 ));
    CascadeMux I__283 (
            .O(N__1882),
            .I(N__1879));
    InMux I__282 (
            .O(N__1879),
            .I(N__1876));
    LocalMux I__281 (
            .O(N__1876),
            .I(\uart_tx.N_143_0 ));
    InMux I__280 (
            .O(N__1873),
            .I(N__1865));
    InMux I__279 (
            .O(N__1872),
            .I(N__1865));
    InMux I__278 (
            .O(N__1871),
            .I(N__1860));
    InMux I__277 (
            .O(N__1870),
            .I(N__1860));
    LocalMux I__276 (
            .O(N__1865),
            .I(\uart_tx.M_bitCtr_qZ0Z_1 ));
    LocalMux I__275 (
            .O(N__1860),
            .I(\uart_tx.M_bitCtr_qZ0Z_1 ));
    CascadeMux I__274 (
            .O(N__1855),
            .I(\uart_tx.M_txReg_q_RNOZ0Z_4_cascade_ ));
    InMux I__273 (
            .O(N__1852),
            .I(N__1849));
    LocalMux I__272 (
            .O(N__1849),
            .I(N__1842));
    InMux I__271 (
            .O(N__1848),
            .I(N__1839));
    InMux I__270 (
            .O(N__1847),
            .I(N__1834));
    InMux I__269 (
            .O(N__1846),
            .I(N__1834));
    InMux I__268 (
            .O(N__1845),
            .I(N__1831));
    Odrv4 I__267 (
            .O(N__1842),
            .I(\uart_tx.M_bitCtr_qZ1Z_0 ));
    LocalMux I__266 (
            .O(N__1839),
            .I(\uart_tx.M_bitCtr_qZ1Z_0 ));
    LocalMux I__265 (
            .O(N__1834),
            .I(\uart_tx.M_bitCtr_qZ1Z_0 ));
    LocalMux I__264 (
            .O(N__1831),
            .I(\uart_tx.M_bitCtr_qZ1Z_0 ));
    InMux I__263 (
            .O(N__1822),
            .I(N__1819));
    LocalMux I__262 (
            .O(N__1819),
            .I(N__1816));
    Odrv4 I__261 (
            .O(N__1816),
            .I(\uart_tx.M_txReg_q_RNOZ0Z_2 ));
    CascadeMux I__260 (
            .O(N__1813),
            .I(\uart_tx.M_txReg_d_3_7_ns_1_cascade_ ));
    InMux I__259 (
            .O(N__1810),
            .I(N__1807));
    LocalMux I__258 (
            .O(N__1807),
            .I(\uart_tx.M_txReg_q_RNOZ0Z_1 ));
    InMux I__257 (
            .O(N__1804),
            .I(N__1796));
    InMux I__256 (
            .O(N__1803),
            .I(N__1785));
    InMux I__255 (
            .O(N__1802),
            .I(N__1785));
    InMux I__254 (
            .O(N__1801),
            .I(N__1785));
    InMux I__253 (
            .O(N__1800),
            .I(N__1785));
    InMux I__252 (
            .O(N__1799),
            .I(N__1785));
    LocalMux I__251 (
            .O(N__1796),
            .I(\uart_tx.M_bitCtr_qZ0Z_2 ));
    LocalMux I__250 (
            .O(N__1785),
            .I(\uart_tx.M_bitCtr_qZ0Z_2 ));
    InMux I__249 (
            .O(N__1780),
            .I(N__1777));
    LocalMux I__248 (
            .O(N__1777),
            .I(\uart_tx.M_txReg_q_RNOZ0Z_5 ));
    InMux I__247 (
            .O(N__1774),
            .I(N__1771));
    LocalMux I__246 (
            .O(N__1771),
            .I(\reset_cond.M_stage_qZ0Z_2 ));
    InMux I__245 (
            .O(N__1768),
            .I(N__1765));
    LocalMux I__244 (
            .O(N__1765),
            .I(N__1759));
    InMux I__243 (
            .O(N__1764),
            .I(N__1752));
    InMux I__242 (
            .O(N__1763),
            .I(N__1752));
    InMux I__241 (
            .O(N__1762),
            .I(N__1752));
    Span4Mux_h I__240 (
            .O(N__1759),
            .I(N__1749));
    LocalMux I__239 (
            .O(N__1752),
            .I(N__1746));
    Sp12to4 I__238 (
            .O(N__1749),
            .I(N__1741));
    Span12Mux_h I__237 (
            .O(N__1746),
            .I(N__1741));
    Span12Mux_v I__236 (
            .O(N__1741),
            .I(N__1738));
    Odrv12 I__235 (
            .O(N__1738),
            .I(rst_n_c));
    InMux I__234 (
            .O(N__1735),
            .I(N__1732));
    LocalMux I__233 (
            .O(N__1732),
            .I(\reset_cond.M_stage_qZ0Z_0 ));
    InMux I__232 (
            .O(N__1729),
            .I(N__1726));
    LocalMux I__231 (
            .O(N__1726),
            .I(\reset_cond.M_stage_qZ0Z_1 ));
    CascadeMux I__230 (
            .O(N__1723),
            .I(N__1719));
    InMux I__229 (
            .O(N__1722),
            .I(N__1716));
    InMux I__228 (
            .O(N__1719),
            .I(N__1713));
    LocalMux I__227 (
            .O(N__1716),
            .I(\uart_tx.N_186_1_i ));
    LocalMux I__226 (
            .O(N__1713),
            .I(\uart_tx.N_186_1_i ));
    InMux I__225 (
            .O(N__1708),
            .I(N__1704));
    InMux I__224 (
            .O(N__1707),
            .I(N__1701));
    LocalMux I__223 (
            .O(N__1704),
            .I(\uart_tx.M_ctr_qZ0Z_0 ));
    LocalMux I__222 (
            .O(N__1701),
            .I(\uart_tx.M_ctr_qZ0Z_0 ));
    CascadeMux I__221 (
            .O(N__1696),
            .I(N__1692));
    InMux I__220 (
            .O(N__1695),
            .I(N__1689));
    InMux I__219 (
            .O(N__1692),
            .I(N__1686));
    LocalMux I__218 (
            .O(N__1689),
            .I(\uart_tx.M_ctr_qZ1Z_1 ));
    LocalMux I__217 (
            .O(N__1686),
            .I(\uart_tx.M_ctr_qZ1Z_1 ));
    InMux I__216 (
            .O(N__1681),
            .I(\uart_tx.un1_M_ctr_q_3_cry_0 ));
    InMux I__215 (
            .O(N__1678),
            .I(N__1674));
    InMux I__214 (
            .O(N__1677),
            .I(N__1671));
    LocalMux I__213 (
            .O(N__1674),
            .I(\uart_tx.M_ctr_qZ0Z_2 ));
    LocalMux I__212 (
            .O(N__1671),
            .I(\uart_tx.M_ctr_qZ0Z_2 ));
    InMux I__211 (
            .O(N__1666),
            .I(N__1663));
    LocalMux I__210 (
            .O(N__1663),
            .I(\uart_tx.M_ctr_q_RNO_0Z0Z_2 ));
    InMux I__209 (
            .O(N__1660),
            .I(\uart_tx.un1_M_ctr_q_3_cry_1 ));
    InMux I__208 (
            .O(N__1657),
            .I(N__1653));
    InMux I__207 (
            .O(N__1656),
            .I(N__1650));
    LocalMux I__206 (
            .O(N__1653),
            .I(\uart_tx.M_ctr_qZ0Z_3 ));
    LocalMux I__205 (
            .O(N__1650),
            .I(\uart_tx.M_ctr_qZ0Z_3 ));
    InMux I__204 (
            .O(N__1645),
            .I(\uart_tx.un1_M_ctr_q_3_cry_2 ));
    InMux I__203 (
            .O(N__1642),
            .I(N__1638));
    InMux I__202 (
            .O(N__1641),
            .I(N__1635));
    LocalMux I__201 (
            .O(N__1638),
            .I(\uart_tx.M_ctr_qZ1Z_4 ));
    LocalMux I__200 (
            .O(N__1635),
            .I(\uart_tx.M_ctr_qZ1Z_4 ));
    InMux I__199 (
            .O(N__1630),
            .I(\uart_tx.un1_M_ctr_q_3_cry_3 ));
    InMux I__198 (
            .O(N__1627),
            .I(N__1623));
    InMux I__197 (
            .O(N__1626),
            .I(N__1620));
    LocalMux I__196 (
            .O(N__1623),
            .I(\uart_tx.M_ctr_qZ1Z_5 ));
    LocalMux I__195 (
            .O(N__1620),
            .I(\uart_tx.M_ctr_qZ1Z_5 ));
    InMux I__194 (
            .O(N__1615),
            .I(N__1612));
    LocalMux I__193 (
            .O(N__1612),
            .I(\uart_tx.M_ctr_q_RNO_0Z0Z_5 ));
    InMux I__192 (
            .O(N__1609),
            .I(\uart_tx.un1_M_ctr_q_3_cry_4 ));
    InMux I__191 (
            .O(N__1606),
            .I(N__1603));
    LocalMux I__190 (
            .O(N__1603),
            .I(un1_M_count_q_axbxc7_1));
    CascadeMux I__189 (
            .O(N__1600),
            .I(\btn_cond.out_17_6_cascade_ ));
    InMux I__188 (
            .O(N__1597),
            .I(N__1594));
    LocalMux I__187 (
            .O(N__1594),
            .I(\btn_cond.out_17_8 ));
    CascadeMux I__186 (
            .O(N__1591),
            .I(btn_cond_out_17_cascade_));
    InMux I__185 (
            .O(N__1588),
            .I(N__1582));
    InMux I__184 (
            .O(N__1587),
            .I(N__1575));
    InMux I__183 (
            .O(N__1586),
            .I(N__1575));
    InMux I__182 (
            .O(N__1585),
            .I(N__1575));
    LocalMux I__181 (
            .O(N__1582),
            .I(N__1572));
    LocalMux I__180 (
            .O(N__1575),
            .I(click_dtct_out8));
    Odrv4 I__179 (
            .O(N__1572),
            .I(click_dtct_out8));
    InMux I__178 (
            .O(N__1567),
            .I(N__1564));
    LocalMux I__177 (
            .O(N__1564),
            .I(\btn_cond.out_17_7 ));
    CascadeMux I__176 (
            .O(N__1561),
            .I(click_dtct_M_count_d6_0_1_cascade_));
    CascadeMux I__175 (
            .O(N__1558),
            .I(\uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_ ));
    InMux I__174 (
            .O(N__1555),
            .I(N__1552));
    LocalMux I__173 (
            .O(N__1552),
            .I(uart_tx_N_187));
    CascadeMux I__172 (
            .O(N__1549),
            .I(un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_));
    InMux I__171 (
            .O(N__1546),
            .I(N__1543));
    LocalMux I__170 (
            .O(N__1543),
            .I(un1_M_count_q_ac0_5_m2_0_a2_3));
    CascadeMux I__169 (
            .O(N__1540),
            .I(un1_M_count_q_ac0_5_m2_0_a2_3_cascade_));
    InMux I__168 (
            .O(N__1537),
            .I(N__1533));
    InMux I__167 (
            .O(N__1536),
            .I(N__1530));
    LocalMux I__166 (
            .O(N__1533),
            .I(un1_M_count_q_ac0_out));
    LocalMux I__165 (
            .O(N__1530),
            .I(un1_M_count_q_ac0_out));
    InMux I__164 (
            .O(N__1525),
            .I(N__1516));
    InMux I__163 (
            .O(N__1524),
            .I(N__1516));
    InMux I__162 (
            .O(N__1523),
            .I(N__1513));
    InMux I__161 (
            .O(N__1522),
            .I(N__1510));
    InMux I__160 (
            .O(N__1521),
            .I(N__1507));
    LocalMux I__159 (
            .O(N__1516),
            .I(click_dtct_out3));
    LocalMux I__158 (
            .O(N__1513),
            .I(click_dtct_out3));
    LocalMux I__157 (
            .O(N__1510),
            .I(click_dtct_out3));
    LocalMux I__156 (
            .O(N__1507),
            .I(click_dtct_out3));
    SRMux I__155 (
            .O(N__1498),
            .I(N__1493));
    SRMux I__154 (
            .O(N__1497),
            .I(N__1490));
    SRMux I__153 (
            .O(N__1496),
            .I(N__1487));
    LocalMux I__152 (
            .O(N__1493),
            .I(N__1484));
    LocalMux I__151 (
            .O(N__1490),
            .I(N__1480));
    LocalMux I__150 (
            .O(N__1487),
            .I(N__1477));
    Span4Mux_v I__149 (
            .O(N__1484),
            .I(N__1474));
    InMux I__148 (
            .O(N__1483),
            .I(N__1471));
    Span4Mux_v I__147 (
            .O(N__1480),
            .I(N__1467));
    Span4Mux_v I__146 (
            .O(N__1477),
            .I(N__1460));
    Span4Mux_h I__145 (
            .O(N__1474),
            .I(N__1460));
    LocalMux I__144 (
            .O(N__1471),
            .I(N__1460));
    InMux I__143 (
            .O(N__1470),
            .I(N__1457));
    Odrv4 I__142 (
            .O(N__1467),
            .I(M_reset_cond_out_0));
    Odrv4 I__141 (
            .O(N__1460),
            .I(M_reset_cond_out_0));
    LocalMux I__140 (
            .O(N__1457),
            .I(M_reset_cond_out_0));
    CascadeMux I__139 (
            .O(N__1450),
            .I(\uart_tx.M_state_q_ns_0_o2_4_0_cascade_ ));
    CascadeMux I__138 (
            .O(N__1447),
            .I(\uart_tx.N_182_0_cascade_ ));
    CascadeMux I__137 (
            .O(N__1444),
            .I(\uart_tx.N_143_0_cascade_ ));
    CascadeMux I__136 (
            .O(N__1441),
            .I(uart_tx_N_185_cascade_));
    InMux I__135 (
            .O(N__1438),
            .I(N__1435));
    LocalMux I__134 (
            .O(N__1435),
            .I(un1_M_count_q_ac0_1));
    CascadeMux I__133 (
            .O(N__1432),
            .I(click_dtct_out3_cascade_));
    CascadeMux I__132 (
            .O(N__1429),
            .I(un1_M_count_q_ac0_7_cascade_));
    InMux I__131 (
            .O(N__1426),
            .I(N__1414));
    InMux I__130 (
            .O(N__1425),
            .I(N__1414));
    InMux I__129 (
            .O(N__1424),
            .I(N__1414));
    InMux I__128 (
            .O(N__1423),
            .I(N__1414));
    LocalMux I__127 (
            .O(N__1414),
            .I(click_dtct_out_d));
    CascadeMux I__126 (
            .O(N__1411),
            .I(click_dtct_out_d_cascade_));
    InMux I__125 (
            .O(N__1408),
            .I(N__1404));
    InMux I__124 (
            .O(N__1407),
            .I(N__1401));
    LocalMux I__123 (
            .O(N__1404),
            .I(un1_M_count_q_ac0_7));
    LocalMux I__122 (
            .O(N__1401),
            .I(un1_M_count_q_ac0_7));
    CascadeMux I__121 (
            .O(N__1396),
            .I(\uart_tx.N_134_i_cascade_ ));
    CascadeMux I__120 (
            .O(N__1393),
            .I(un1_M_count_q_ac0_1_cascade_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(\btn_cond.un1_M_ctr_q_cry_7 ),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(\btn_cond.un1_M_ctr_q_cry_15 ),
            .carryinitout(bfn_15_27_0_));
    ICE_GB \btn_cond.sync.M_pipe_q_RNIJLM5_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__2842),
            .GLOBALBUFFEROUTPUT(\btn_cond.M_sync_out_i_g_0 ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam M_count_q_RNI2B741_0_LC_13_23_3.C_ON=1'b0;
    defparam M_count_q_RNI2B741_0_LC_13_23_3.SEQ_MODE=4'b0000;
    defparam M_count_q_RNI2B741_0_LC_13_23_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 M_count_q_RNI2B741_0_LC_13_23_3 (
            .in0(_gnd_net_),
            .in1(N__2234),
            .in2(_gnd_net_),
            .in3(N__2303),
            .lcout(un1_M_count_q_ac0_out),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNI0H5P2_1_LC_13_24_0.C_ON=1'b0;
    defparam M_count_q_RNI0H5P2_1_LC_13_24_0.SEQ_MODE=4'b0000;
    defparam M_count_q_RNI0H5P2_1_LC_13_24_0.LUT_INIT=16'b1000100010000000;
    LogicCell40 M_count_q_RNI0H5P2_1_LC_13_24_0 (
            .in0(N__2765),
            .in1(N__1536),
            .in2(N__2008),
            .in3(N__1521),
            .lcout(un1_M_count_q_ac0_1),
            .ltout(un1_M_count_q_ac0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_2_LC_13_24_1.C_ON=1'b0;
    defparam M_count_q_2_LC_13_24_1.SEQ_MODE=4'b1000;
    defparam M_count_q_2_LC_13_24_1.LUT_INIT=16'b0011110011001100;
    LogicCell40 M_count_q_2_LC_13_24_1 (
            .in0(_gnd_net_),
            .in1(N__2819),
            .in2(N__1393),
            .in3(N__1423),
            .lcout(M_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2900),
            .ce(),
            .sr(N__1498));
    defparam M_count_q_5_LC_13_24_3.C_ON=1'b0;
    defparam M_count_q_5_LC_13_24_3.SEQ_MODE=4'b1000;
    defparam M_count_q_5_LC_13_24_3.LUT_INIT=16'b0110011010101010;
    LogicCell40 M_count_q_5_LC_13_24_3 (
            .in0(N__2723),
            .in1(N__1424),
            .in2(_gnd_net_),
            .in3(N__1407),
            .lcout(M_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2900),
            .ce(),
            .sr(N__1498));
    defparam M_count_q_3_LC_13_24_4.C_ON=1'b0;
    defparam M_count_q_3_LC_13_24_4.SEQ_MODE=4'b1000;
    defparam M_count_q_3_LC_13_24_4.LUT_INIT=16'b0110110011001100;
    LogicCell40 M_count_q_3_LC_13_24_4 (
            .in0(N__1425),
            .in1(N__2790),
            .in2(N__2826),
            .in3(N__1438),
            .lcout(M_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2900),
            .ce(),
            .sr(N__1498));
    defparam \click_dtct.M_last_q_RNIUTK51_1_LC_13_24_5 .C_ON=1'b0;
    defparam \click_dtct.M_last_q_RNIUTK51_1_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \click_dtct.M_last_q_RNIUTK51_1_LC_13_24_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \click_dtct.M_last_q_RNIUTK51_1_LC_13_24_5  (
            .in0(N__2088),
            .in1(N__2064),
            .in2(N__2006),
            .in3(N__2029),
            .lcout(click_dtct_out3),
            .ltout(click_dtct_out3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIGFD24_4_LC_13_24_6.C_ON=1'b0;
    defparam M_count_q_RNIGFD24_4_LC_13_24_6.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIGFD24_4_LC_13_24_6.LUT_INIT=16'b1000100010000000;
    LogicCell40 M_count_q_RNIGFD24_4_LC_13_24_6 (
            .in0(N__1546),
            .in1(N__2162),
            .in2(N__1432),
            .in3(N__1997),
            .lcout(un1_M_count_q_ac0_7),
            .ltout(un1_M_count_q_ac0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_6_LC_13_24_7.C_ON=1'b0;
    defparam M_count_q_6_LC_13_24_7.SEQ_MODE=4'b1000;
    defparam M_count_q_6_LC_13_24_7.LUT_INIT=16'b0110110011001100;
    LogicCell40 M_count_q_6_LC_13_24_7 (
            .in0(N__2724),
            .in1(N__2199),
            .in2(N__1429),
            .in3(N__1426),
            .lcout(M_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2900),
            .ce(),
            .sr(N__1498));
    defparam \click_dtct.M_last_q_RNIUTK51_LC_13_25_1 .C_ON=1'b0;
    defparam \click_dtct.M_last_q_RNIUTK51_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \click_dtct.M_last_q_RNIUTK51_LC_13_25_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \click_dtct.M_last_q_RNIUTK51_LC_13_25_1  (
            .in0(N__2090),
            .in1(N__2061),
            .in2(N__2007),
            .in3(N__2031),
            .lcout(click_dtct_out_d),
            .ltout(click_dtct_out_d_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_7_LC_13_25_2.C_ON=1'b0;
    defparam M_count_q_7_LC_13_25_2.SEQ_MODE=4'b1000;
    defparam M_count_q_7_LC_13_25_2.LUT_INIT=16'b1001101010101010;
    LogicCell40 M_count_q_7_LC_13_25_2 (
            .in0(N__2133),
            .in1(N__1606),
            .in2(N__1411),
            .in3(N__1408),
            .lcout(M_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2903),
            .ce(),
            .sr(N__1496));
    defparam \reset_cond.M_stage_q_3_LC_14_21_0 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_3_LC_14_21_0 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_3_LC_14_21_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \reset_cond.M_stage_q_3_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__1768),
            .in2(_gnd_net_),
            .in3(N__1774),
            .lcout(M_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2892),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_5_LC_14_22_0 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_5_LC_14_22_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_5_LC_14_22_0 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \uart_tx.M_ctr_q_5_LC_14_22_0  (
            .in0(N__2313),
            .in1(N__1615),
            .in2(N__1942),
            .in3(N__1922),
            .lcout(\uart_tx.M_ctr_qZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2895),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_RNILEFM_0_1_LC_14_22_1 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNILEFM_0_1_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNILEFM_0_1_LC_14_22_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uart_tx.M_state_q_RNILEFM_0_1_LC_14_22_1  (
            .in0(N__2377),
            .in1(_gnd_net_),
            .in2(N__2435),
            .in3(_gnd_net_),
            .lcout(\uart_tx.N_134_i ),
            .ltout(\uart_tx.N_134_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_2_LC_14_22_2 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_2_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_2_LC_14_22_2 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \uart_tx.M_ctr_q_2_LC_14_22_2  (
            .in0(N__2312),
            .in1(N__1666),
            .in2(N__1396),
            .in3(N__1921),
            .lcout(\uart_tx.M_ctr_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2895),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_1_LC_14_22_3 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_1_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_state_q_1_LC_14_22_3 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \uart_tx.M_state_q_1_LC_14_22_3  (
            .in0(N__1923),
            .in1(N__1470),
            .in2(N__2388),
            .in3(N__2434),
            .lcout(\uart_tx.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2895),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_RNILEFM_1_LC_14_22_4 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNILEFM_1_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNILEFM_1_LC_14_22_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_tx.M_state_q_RNILEFM_1_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__2420),
            .in2(_gnd_net_),
            .in3(N__2376),
            .lcout(\uart_tx.N_186_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNIGGUF1_0_LC_14_22_5 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_RNIGGUF1_0_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNIGGUF1_0_LC_14_22_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uart_tx.M_ctr_q_RNIGGUF1_0_LC_14_22_5  (
            .in0(N__1626),
            .in1(N__1677),
            .in2(N__1696),
            .in3(N__1707),
            .lcout(),
            .ltout(\uart_tx.M_state_q_ns_0_o2_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNI3KTJ2_6_LC_14_22_6 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_RNI3KTJ2_6_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNI3KTJ2_6_LC_14_22_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_tx.M_ctr_q_RNI3KTJ2_6_LC_14_22_6  (
            .in0(N__1893),
            .in1(N__1641),
            .in2(N__1450),
            .in3(N__1656),
            .lcout(\uart_tx.N_182_0 ),
            .ltout(\uart_tx.N_182_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_0_LC_14_22_7 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_0_LC_14_22_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_bitCtr_q_0_LC_14_22_7 .LUT_INIT=16'b1100110000101000;
    LogicCell40 \uart_tx.M_bitCtr_q_0_LC_14_22_7  (
            .in0(N__2378),
            .in1(N__1852),
            .in2(N__1447),
            .in3(N__2433),
            .lcout(\uart_tx.M_bitCtr_qZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2895),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_RNIP5AF3_0_LC_14_23_0 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_RNIP5AF3_0_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_bitCtr_q_RNIP5AF3_0_LC_14_23_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uart_tx.M_bitCtr_q_RNIP5AF3_0_LC_14_23_0  (
            .in0(N__2384),
            .in1(N__1848),
            .in2(N__2436),
            .in3(N__1920),
            .lcout(\uart_tx.N_143_0 ),
            .ltout(\uart_tx.N_143_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_1_LC_14_23_1 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_1_LC_14_23_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_bitCtr_q_1_LC_14_23_1 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \uart_tx.M_bitCtr_q_1_LC_14_23_1  (
            .in0(N__1871),
            .in1(_gnd_net_),
            .in2(N__1444),
            .in3(N__2311),
            .lcout(\uart_tx.M_bitCtr_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2897),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_RNITA5V2_0_LC_14_23_2 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNITA5V2_0_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNITA5V2_0_LC_14_23_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uart_tx.M_state_q_RNITA5V2_0_LC_14_23_2  (
            .in0(N__2426),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1918),
            .lcout(),
            .ltout(uart_tx_N_185_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \click_dtct.M_last_q_RNIE6EK8_LC_14_23_3 .C_ON=1'b0;
    defparam \click_dtct.M_last_q_RNIE6EK8_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \click_dtct.M_last_q_RNIE6EK8_LC_14_23_3 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \click_dtct.M_last_q_RNIE6EK8_LC_14_23_3  (
            .in0(N__1522),
            .in1(N__2309),
            .in2(N__1441),
            .in3(N__1555),
            .lcout(),
            .ltout(click_dtct_M_count_d6_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_0_LC_14_23_4 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_0_LC_14_23_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_state_q_0_LC_14_23_4 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \uart_tx.M_state_q_0_LC_14_23_4  (
            .in0(N__2310),
            .in1(N__1483),
            .in2(N__1561),
            .in3(N__1588),
            .lcout(\uart_tx.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2897),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_RNITT1L_1_LC_14_23_5 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_RNITT1L_1_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_bitCtr_q_RNITT1L_1_LC_14_23_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_tx.M_bitCtr_q_RNITT1L_1_LC_14_23_5  (
            .in0(N__1870),
            .in1(N__1845),
            .in2(_gnd_net_),
            .in3(N__2425),
            .lcout(),
            .ltout(\uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_RNIUE4P3_2_LC_14_23_6 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_RNIUE4P3_2_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_bitCtr_q_RNIUE4P3_2_LC_14_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_tx.M_bitCtr_q_RNIUE4P3_2_LC_14_23_6  (
            .in0(N__2383),
            .in1(N__1804),
            .in2(N__1558),
            .in3(N__1919),
            .lcout(uart_tx_N_187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_RNILEFM_1_1_LC_14_23_7 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNILEFM_1_1_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNILEFM_1_1_LC_14_23_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_tx.M_state_q_RNILEFM_1_1_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__2424),
            .in2(_gnd_net_),
            .in3(N__2382),
            .lcout(uart_tx_N_186_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_0_LC_14_24_1.C_ON=1'b0;
    defparam M_count_q_0_LC_14_24_1.SEQ_MODE=4'b1000;
    defparam M_count_q_0_LC_14_24_1.LUT_INIT=16'b0101101001111000;
    LogicCell40 M_count_q_0_LC_14_24_1 (
            .in0(N__2317),
            .in1(N__1585),
            .in2(N__2238),
            .in3(N__1524),
            .lcout(M_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2898),
            .ce(),
            .sr(N__1497));
    defparam M_count_q_RNITRFR_3_LC_14_24_2.C_ON=1'b0;
    defparam M_count_q_RNITRFR_3_LC_14_24_2.SEQ_MODE=4'b0000;
    defparam M_count_q_RNITRFR_3_LC_14_24_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 M_count_q_RNITRFR_3_LC_14_24_2 (
            .in0(_gnd_net_),
            .in1(N__2789),
            .in2(_gnd_net_),
            .in3(N__2230),
            .lcout(),
            .ltout(un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIF6FD2_1_LC_14_24_3.C_ON=1'b0;
    defparam M_count_q_RNIF6FD2_1_LC_14_24_3.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIF6FD2_1_LC_14_24_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_count_q_RNIF6FD2_1_LC_14_24_3 (
            .in0(N__2818),
            .in1(N__2755),
            .in2(N__1549),
            .in3(N__2304),
            .lcout(un1_M_count_q_ac0_5_m2_0_a2_3),
            .ltout(un1_M_count_q_ac0_5_m2_0_a2_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_4_LC_14_24_4.C_ON=1'b0;
    defparam M_count_q_4_LC_14_24_4.SEQ_MODE=4'b1000;
    defparam M_count_q_4_LC_14_24_4.LUT_INIT=16'b0001111111100000;
    LogicCell40 M_count_q_4_LC_14_24_4 (
            .in0(N__1587),
            .in1(N__1523),
            .in2(N__1540),
            .in3(N__2163),
            .lcout(M_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2898),
            .ce(),
            .sr(N__1497));
    defparam M_count_q_1_LC_14_24_5.C_ON=1'b0;
    defparam M_count_q_1_LC_14_24_5.SEQ_MODE=4'b1000;
    defparam M_count_q_1_LC_14_24_5.LUT_INIT=16'b0101101001111000;
    LogicCell40 M_count_q_1_LC_14_24_5 (
            .in0(N__1537),
            .in1(N__1586),
            .in2(N__2766),
            .in3(N__1525),
            .lcout(M_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2898),
            .ce(),
            .sr(N__1497));
    defparam \btn_cond.M_ctr_q_RNIUMNB_4_LC_14_25_1 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIUMNB_4_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIUMNB_4_LC_14_25_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \btn_cond.M_ctr_q_RNIUMNB_4_LC_14_25_1  (
            .in0(N__2664),
            .in1(N__2682),
            .in2(N__2626),
            .in3(N__2645),
            .lcout(\btn_cond.out_17_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNO_0_7_LC_14_25_2.C_ON=1'b0;
    defparam M_count_q_RNO_0_7_LC_14_25_2.SEQ_MODE=4'b0000;
    defparam M_count_q_RNO_0_7_LC_14_25_2.LUT_INIT=16'b0101010111111111;
    LogicCell40 M_count_q_RNO_0_7_LC_14_25_2 (
            .in0(N__2714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2198),
            .lcout(un1_M_count_q_axbxc7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIE6NB_0_LC_14_25_3 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIE6NB_0_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIE6NB_0_LC_14_25_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \btn_cond.M_ctr_q_RNIE6NB_0_LC_14_25_3  (
            .in0(N__3096),
            .in1(N__3158),
            .in2(N__3121),
            .in3(N__3138),
            .lcout(btn_cond_out_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIQGM2_12_LC_14_25_4 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIQGM2_12_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIQGM2_12_LC_14_25_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \btn_cond.M_ctr_q_RNIQGM2_12_LC_14_25_4  (
            .in0(N__3055),
            .in1(N__3072),
            .in2(N__2521),
            .in3(N__2498),
            .lcout(),
            .ltout(\btn_cond.out_17_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIKBLL_10_LC_14_25_5 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIKBLL_10_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIKBLL_10_LC_14_25_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \btn_cond.M_ctr_q_RNIKBLL_10_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__1567),
            .in2(N__1600),
            .in3(N__1597),
            .lcout(btn_cond_out_17),
            .ltout(btn_cond_out_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \click_dtct.M_last_q_RNIUTK51_0_LC_14_25_6 .C_ON=1'b0;
    defparam \click_dtct.M_last_q_RNIUTK51_0_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \click_dtct.M_last_q_RNIUTK51_0_LC_14_25_6 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \click_dtct.M_last_q_RNIUTK51_0_LC_14_25_6  (
            .in0(N__2004),
            .in1(N__2062),
            .in2(N__1591),
            .in3(N__2091),
            .lcout(click_dtct_out8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \click_dtct.M_last_q_LC_14_25_7 .C_ON=1'b0;
    defparam \click_dtct.M_last_q_LC_14_25_7 .SEQ_MODE=4'b1000;
    defparam \click_dtct.M_last_q_LC_14_25_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \click_dtct.M_last_q_LC_14_25_7  (
            .in0(N__2063),
            .in1(_gnd_net_),
            .in2(N__2095),
            .in3(N__2032),
            .lcout(click_dtct_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2901),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIA1N2_19_LC_14_26_1 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIA1N2_19_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIA1N2_19_LC_14_26_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \btn_cond.M_ctr_q_RNIA1N2_19_LC_14_26_1  (
            .in0(N__3007),
            .in1(N__2984),
            .in2(N__2965),
            .in3(N__3024),
            .lcout(btn_cond_out_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIS377_10_LC_14_26_4 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIS377_10_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIS377_10_LC_14_26_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \btn_cond.M_ctr_q_RNIS377_10_LC_14_26_4  (
            .in0(N__2602),
            .in1(N__2558),
            .in2(N__2581),
            .in3(N__2538),
            .lcout(\btn_cond.out_17_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_0_LC_15_21_3 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_0_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_0_LC_15_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \reset_cond.M_stage_q_0_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1762),
            .lcout(\reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2890),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_2_LC_15_21_4 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_2_LC_15_21_4 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_2_LC_15_21_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \reset_cond.M_stage_q_2_LC_15_21_4  (
            .in0(N__1764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1729),
            .lcout(\reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2890),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_1_LC_15_21_5 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_1_LC_15_21_5 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_1_LC_15_21_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \reset_cond.M_stage_q_1_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__1763),
            .in2(_gnd_net_),
            .in3(N__1735),
            .lcout(\reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2890),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_0_LC_15_22_0 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_0_LC_15_22_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_0_LC_15_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_0_LC_15_22_0  (
            .in0(N__2314),
            .in1(N__1708),
            .in2(N__1723),
            .in3(N__1722),
            .lcout(\uart_tx.M_ctr_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_0 ),
            .clk(N__2893),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_1_LC_15_22_1 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_1_LC_15_22_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_1_LC_15_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_1_LC_15_22_1  (
            .in0(N__2327),
            .in1(N__1695),
            .in2(_gnd_net_),
            .in3(N__1681),
            .lcout(\uart_tx.M_ctr_qZ1Z_1 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_0 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_1 ),
            .clk(N__2893),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNO_0_2_LC_15_22_2 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_RNO_0_2_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNO_0_2_LC_15_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.M_ctr_q_RNO_0_2_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__1678),
            .in2(_gnd_net_),
            .in3(N__1660),
            .lcout(\uart_tx.M_ctr_q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_1 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_3_LC_15_22_3 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_3_LC_15_22_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_3_LC_15_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_3_LC_15_22_3  (
            .in0(N__2328),
            .in1(N__1657),
            .in2(_gnd_net_),
            .in3(N__1645),
            .lcout(\uart_tx.M_ctr_qZ0Z_3 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_2 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_3 ),
            .clk(N__2893),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_4_LC_15_22_4 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_4_LC_15_22_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_4_LC_15_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_4_LC_15_22_4  (
            .in0(N__2315),
            .in1(N__1642),
            .in2(_gnd_net_),
            .in3(N__1630),
            .lcout(\uart_tx.M_ctr_qZ1Z_4 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_3 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_4 ),
            .clk(N__2893),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNO_0_5_LC_15_22_5 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_RNO_0_5_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNO_0_5_LC_15_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.M_ctr_q_RNO_0_5_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__1627),
            .in2(_gnd_net_),
            .in3(N__1609),
            .lcout(\uart_tx.M_ctr_q_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_4 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNO_0_6_LC_15_22_6 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_RNO_0_6_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNO_0_6_LC_15_22_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_tx.M_ctr_q_RNO_0_6_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__1894),
            .in2(_gnd_net_),
            .in3(N__1945),
            .lcout(),
            .ltout(\uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_6_LC_15_22_7 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_6_LC_15_22_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_6_LC_15_22_7 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \uart_tx.M_ctr_q_6_LC_15_22_7  (
            .in0(N__1941),
            .in1(N__2316),
            .in2(N__1927),
            .in3(N__1924),
            .lcout(\uart_tx.M_ctr_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2893),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_2_LC_15_23_0 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_2_LC_15_23_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_bitCtr_q_2_LC_15_23_0 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uart_tx.M_bitCtr_q_2_LC_15_23_0  (
            .in0(N__1803),
            .in1(N__1873),
            .in2(N__1882),
            .in3(N__2323),
            .lcout(\uart_tx.M_bitCtr_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2896),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_2_LC_15_23_1 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_2_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_2_LC_15_23_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uart_tx.M_txReg_q_RNO_2_LC_15_23_1  (
            .in0(N__2773),
            .in1(N__2836),
            .in2(_gnd_net_),
            .in3(N__1802),
            .lcout(\uart_tx.M_txReg_q_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_4_LC_15_23_2 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_4_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_4_LC_15_23_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart_tx.M_txReg_q_RNO_4_LC_15_23_2  (
            .in0(N__1800),
            .in1(N__2146),
            .in2(_gnd_net_),
            .in3(N__2212),
            .lcout(),
            .ltout(\uart_tx.M_txReg_q_RNOZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_3_LC_15_23_3 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_3_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_3_LC_15_23_3 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \uart_tx.M_txReg_q_RNO_3_LC_15_23_3  (
            .in0(N__1872),
            .in1(N__1846),
            .in2(N__1855),
            .in3(N__1780),
            .lcout(),
            .ltout(\uart_tx.M_txReg_d_3_7_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_0_LC_15_23_4 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_0_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_0_LC_15_23_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \uart_tx.M_txReg_q_RNO_0_LC_15_23_4  (
            .in0(N__1847),
            .in1(N__1822),
            .in2(N__1813),
            .in3(N__1810),
            .lcout(\uart_tx.M_txReg_d_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_1_LC_15_23_6 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_1_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_1_LC_15_23_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart_tx.M_txReg_q_RNO_1_LC_15_23_6  (
            .in0(N__1801),
            .in1(N__2701),
            .in2(_gnd_net_),
            .in3(N__2734),
            .lcout(\uart_tx.M_txReg_q_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_5_LC_15_23_7 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_5_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_5_LC_15_23_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uart_tx.M_txReg_q_RNO_5_LC_15_23_7  (
            .in0(N__2800),
            .in1(N__2176),
            .in2(_gnd_net_),
            .in3(N__1799),
            .lcout(\uart_tx.M_txReg_q_RNOZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNICJ341_19_LC_15_24_1 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNICJ341_19_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNICJ341_19_LC_15_24_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \btn_cond.M_ctr_q_RNICJ341_19_LC_15_24_1  (
            .in0(N__2089),
            .in1(N__2065),
            .in2(_gnd_net_),
            .in3(N__2030),
            .lcout(),
            .ltout(M_btn_cond_out_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \click_dtct.M_last_q_RNIJC4S1_LC_15_24_2 .C_ON=1'b0;
    defparam \click_dtct.M_last_q_RNIJC4S1_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \click_dtct.M_last_q_RNIJC4S1_LC_15_24_2 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \click_dtct.M_last_q_RNIJC4S1_LC_15_24_2  (
            .in0(N__2005),
            .in1(_gnd_net_),
            .in2(N__1966),
            .in3(N__2305),
            .lcout(M_count_d6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_0_LC_15_25_0 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_0_LC_15_25_0 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_0_LC_15_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_0_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__3139),
            .in2(N__3175),
            .in3(N__3174),
            .lcout(\btn_cond.M_ctr_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(\btn_cond.un1_M_ctr_q_cry_0 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_1_LC_15_25_1 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_1_LC_15_25_1 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_1_LC_15_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_1_LC_15_25_1  (
            .in0(_gnd_net_),
            .in1(N__3097),
            .in2(_gnd_net_),
            .in3(N__1963),
            .lcout(\btn_cond.M_ctr_qZ0Z_1 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_0 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_1 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_2_LC_15_25_2 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_2_LC_15_25_2 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_2_LC_15_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_2_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__3159),
            .in2(_gnd_net_),
            .in3(N__1960),
            .lcout(\btn_cond.M_ctr_qZ0Z_2 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_1 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_2 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_3_LC_15_25_3 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_3_LC_15_25_3 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_3_LC_15_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_3_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(N__3119),
            .in2(_gnd_net_),
            .in3(N__1957),
            .lcout(\btn_cond.M_ctr_qZ0Z_3 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_2 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_3 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_4_LC_15_25_4 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_4_LC_15_25_4 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_4_LC_15_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_4_LC_15_25_4  (
            .in0(_gnd_net_),
            .in1(N__2646),
            .in2(_gnd_net_),
            .in3(N__1954),
            .lcout(\btn_cond.M_ctr_qZ0Z_4 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_3 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_4 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_5_LC_15_25_5 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_5_LC_15_25_5 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_5_LC_15_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_5_LC_15_25_5  (
            .in0(_gnd_net_),
            .in1(N__2665),
            .in2(_gnd_net_),
            .in3(N__1951),
            .lcout(\btn_cond.M_ctr_qZ0Z_5 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_4 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_5 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_6_LC_15_25_6 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_6_LC_15_25_6 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_6_LC_15_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_6_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(N__2683),
            .in2(_gnd_net_),
            .in3(N__1948),
            .lcout(\btn_cond.M_ctr_qZ0Z_6 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_5 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_6 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_7_LC_15_25_7 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_7_LC_15_25_7 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_7_LC_15_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_7_LC_15_25_7  (
            .in0(_gnd_net_),
            .in1(N__2622),
            .in2(_gnd_net_),
            .in3(N__2122),
            .lcout(\btn_cond.M_ctr_qZ0Z_7 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_6 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_7 ),
            .clk(N__2899),
            .ce(),
            .sr(N__2461));
    defparam \btn_cond.M_ctr_q_8_LC_15_26_0 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_8_LC_15_26_0 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_8_LC_15_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_8_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(N__2580),
            .in2(_gnd_net_),
            .in3(N__2119),
            .lcout(\btn_cond.M_ctr_qZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(\btn_cond.un1_M_ctr_q_cry_8 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_9_LC_15_26_1 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_9_LC_15_26_1 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_9_LC_15_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_9_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__2539),
            .in2(_gnd_net_),
            .in3(N__2116),
            .lcout(\btn_cond.M_ctr_qZ0Z_9 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_8 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_9 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_10_LC_15_26_2 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_10_LC_15_26_2 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_10_LC_15_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_10_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__2559),
            .in2(_gnd_net_),
            .in3(N__2113),
            .lcout(\btn_cond.M_ctr_qZ0Z_10 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_9 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_10 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_11_LC_15_26_3 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_11_LC_15_26_3 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_11_LC_15_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_11_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(N__2601),
            .in2(_gnd_net_),
            .in3(N__2110),
            .lcout(\btn_cond.M_ctr_qZ0Z_11 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_10 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_11 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_12_LC_15_26_4 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_12_LC_15_26_4 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_12_LC_15_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_12_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(N__3073),
            .in2(_gnd_net_),
            .in3(N__2107),
            .lcout(\btn_cond.M_ctr_qZ0Z_12 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_11 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_12 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_13_LC_15_26_5 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_13_LC_15_26_5 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_13_LC_15_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_13_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(N__3051),
            .in2(_gnd_net_),
            .in3(N__2104),
            .lcout(\btn_cond.M_ctr_qZ0Z_13 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_12 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_13 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_14_LC_15_26_6 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_14_LC_15_26_6 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_14_LC_15_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_14_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(N__2500),
            .in2(_gnd_net_),
            .in3(N__2101),
            .lcout(\btn_cond.M_ctr_qZ0Z_14 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_13 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_14 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_15_LC_15_26_7 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_15_LC_15_26_7 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_15_LC_15_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_15_LC_15_26_7  (
            .in0(_gnd_net_),
            .in1(N__2520),
            .in2(_gnd_net_),
            .in3(N__2098),
            .lcout(\btn_cond.M_ctr_qZ0Z_15 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_14 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_15 ),
            .clk(N__2902),
            .ce(),
            .sr(N__2460));
    defparam \btn_cond.M_ctr_q_16_LC_15_27_0 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_16_LC_15_27_0 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_16_LC_15_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_16_LC_15_27_0  (
            .in0(_gnd_net_),
            .in1(N__2961),
            .in2(_gnd_net_),
            .in3(N__2473),
            .lcout(\btn_cond.M_ctr_qZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(\btn_cond.un1_M_ctr_q_cry_16 ),
            .clk(N__2904),
            .ce(),
            .sr(N__2459));
    defparam \btn_cond.M_ctr_q_17_LC_15_27_1 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_17_LC_15_27_1 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_17_LC_15_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_17_LC_15_27_1  (
            .in0(_gnd_net_),
            .in1(N__3006),
            .in2(_gnd_net_),
            .in3(N__2470),
            .lcout(\btn_cond.M_ctr_qZ0Z_17 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_16 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_17 ),
            .clk(N__2904),
            .ce(),
            .sr(N__2459));
    defparam \btn_cond.M_ctr_q_18_LC_15_27_2 .C_ON=1'b1;
    defparam \btn_cond.M_ctr_q_18_LC_15_27_2 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_18_LC_15_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \btn_cond.M_ctr_q_18_LC_15_27_2  (
            .in0(_gnd_net_),
            .in1(N__3025),
            .in2(_gnd_net_),
            .in3(N__2467),
            .lcout(\btn_cond.M_ctr_qZ0Z_18 ),
            .ltout(),
            .carryin(\btn_cond.un1_M_ctr_q_cry_17 ),
            .carryout(\btn_cond.un1_M_ctr_q_cry_18 ),
            .clk(N__2904),
            .ce(),
            .sr(N__2459));
    defparam \btn_cond.M_ctr_q_19_LC_15_27_3 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_19_LC_15_27_3 .SEQ_MODE=4'b1000;
    defparam \btn_cond.M_ctr_q_19_LC_15_27_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \btn_cond.M_ctr_q_19_LC_15_27_3  (
            .in0(_gnd_net_),
            .in1(N__2985),
            .in2(_gnd_net_),
            .in3(N__2464),
            .lcout(\btn_cond.M_ctr_qZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2904),
            .ce(),
            .sr(N__2459));
    defparam \uart_tx.M_txReg_q_LC_16_22_3 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_LC_16_22_3 .SEQ_MODE=4'b1001;
    defparam \uart_tx.M_txReg_q_LC_16_22_3 .LUT_INIT=16'b1110111000110011;
    LogicCell40 \uart_tx.M_txReg_q_LC_16_22_3  (
            .in0(N__2446),
            .in1(N__2440),
            .in2(_gnd_net_),
            .in3(N__2389),
            .lcout(usb_tx_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2889),
            .ce(),
            .sr(N__2329));
    defparam \uart_tx.M_savedData_q_0_LC_16_23_0 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_0_LC_16_23_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_0_LC_16_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_0_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2242),
            .lcout(\uart_tx.M_savedData_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2891),
            .ce(N__2695),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_6_LC_16_23_1 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_6_LC_16_23_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_6_LC_16_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_6_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2203),
            .lcout(\uart_tx.M_savedData_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2891),
            .ce(N__2695),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_4_LC_16_23_4 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_4_LC_16_23_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_4_LC_16_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_4_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2170),
            .lcout(\uart_tx.M_savedData_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2891),
            .ce(N__2695),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_7_LC_16_23_7 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_7_LC_16_23_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_7_LC_16_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_7_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2140),
            .lcout(\uart_tx.M_savedData_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2891),
            .ce(N__2695),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_2_LC_16_24_0 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_2_LC_16_24_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_2_LC_16_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_2_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2827),
            .lcout(\uart_tx.M_savedData_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2894),
            .ce(N__2694),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_3_LC_16_24_1 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_3_LC_16_24_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_3_LC_16_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_3_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2794),
            .lcout(\uart_tx.M_savedData_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2894),
            .ce(N__2694),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_1_LC_16_24_3 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_1_LC_16_24_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_1_LC_16_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_1_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2767),
            .lcout(\uart_tx.M_savedData_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2894),
            .ce(N__2694),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_5_LC_16_24_7 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_5_LC_16_24_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_5_LC_16_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.M_savedData_q_5_LC_16_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2728),
            .lcout(\uart_tx.M_savedData_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2894),
            .ce(N__2694),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIUMNB_0_4_LC_16_25_0 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIUMNB_0_4_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIUMNB_0_4_LC_16_25_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \btn_cond.M_ctr_q_RNIUMNB_0_4_LC_16_25_0  (
            .in0(N__2681),
            .in1(N__2663),
            .in2(N__2647),
            .in3(N__2618),
            .lcout(\btn_cond.g0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIS377_0_10_LC_16_25_2 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIS377_0_10_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIS377_0_10_LC_16_25_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \btn_cond.M_ctr_q_RNIS377_0_10_LC_16_25_2  (
            .in0(N__2597),
            .in1(N__2576),
            .in2(N__2560),
            .in3(N__2537),
            .lcout(),
            .ltout(\btn_cond.g0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIMKT9_14_LC_16_25_3 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIMKT9_14_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIMKT9_14_LC_16_25_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \btn_cond.M_ctr_q_RNIMKT9_14_LC_16_25_3  (
            .in0(N__2516),
            .in1(N__2499),
            .in2(N__2482),
            .in3(N__3031),
            .lcout(),
            .ltout(\btn_cond.g0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNICJ341_14_LC_16_25_4 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNICJ341_14_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNICJ341_14_LC_16_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \btn_cond.M_ctr_q_RNICJ341_14_LC_16_25_4  (
            .in0(N__2479),
            .in1(N__3079),
            .in2(N__3178),
            .in3(N__2941),
            .lcout(\btn_cond.M_btn_cond_out_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIE6NB_0_0_LC_16_25_5 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIE6NB_0_0_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIE6NB_0_0_LC_16_25_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \btn_cond.M_ctr_q_RNIE6NB_0_0_LC_16_25_5  (
            .in0(N__3160),
            .in1(N__3137),
            .in2(N__3120),
            .in3(N__3095),
            .lcout(\btn_cond.g0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIB6B1_12_LC_16_25_7 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIB6B1_12_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIB6B1_12_LC_16_25_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \btn_cond.M_ctr_q_RNIB6B1_12_LC_16_25_7  (
            .in0(_gnd_net_),
            .in1(N__3071),
            .in2(_gnd_net_),
            .in3(N__3047),
            .lcout(\btn_cond.g0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.M_ctr_q_RNIA1N2_0_19_LC_16_26_2 .C_ON=1'b0;
    defparam \btn_cond.M_ctr_q_RNIA1N2_0_19_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \btn_cond.M_ctr_q_RNIA1N2_0_19_LC_16_26_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \btn_cond.M_ctr_q_RNIA1N2_0_19_LC_16_26_2  (
            .in0(N__3023),
            .in1(N__3002),
            .in2(N__2986),
            .in3(N__2957),
            .lcout(\btn_cond.g0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.sync.M_pipe_q_1_LC_16_31_4 .C_ON=1'b0;
    defparam \btn_cond.sync.M_pipe_q_1_LC_16_31_4 .SEQ_MODE=4'b1000;
    defparam \btn_cond.sync.M_pipe_q_1_LC_16_31_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \btn_cond.sync.M_pipe_q_1_LC_16_31_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2911),
            .lcout(\btn_cond.sync.M_sync_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2905),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.sync.M_pipe_q_0_LC_16_31_5 .C_ON=1'b0;
    defparam \btn_cond.sync.M_pipe_q_0_LC_16_31_5 .SEQ_MODE=4'b1000;
    defparam \btn_cond.sync.M_pipe_q_0_LC_16_31_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \btn_cond.sync.M_pipe_q_0_LC_16_31_5  (
            .in0(N__2935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\btn_cond.sync.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2905),
            .ce(),
            .sr(_gnd_net_));
    defparam \btn_cond.sync.M_pipe_q_RNIJLM5_1_LC_16_32_6 .C_ON=1'b0;
    defparam \btn_cond.sync.M_pipe_q_RNIJLM5_1_LC_16_32_6 .SEQ_MODE=4'b0000;
    defparam \btn_cond.sync.M_pipe_q_RNIJLM5_1_LC_16_32_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \btn_cond.sync.M_pipe_q_RNIJLM5_1_LC_16_32_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2848),
            .lcout(\btn_cond.sync.M_sync_out_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
