// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     Oct 30 2022 12:29:41

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    sr_latch,
    sr_data,
    sr_clk,
    rst_n,
    clk);

    output sr_latch;
    output sr_data;
    output sr_clk;
    input rst_n;
    input clk;

    wire N__5116;
    wire N__5115;
    wire N__5114;
    wire N__5105;
    wire N__5104;
    wire N__5103;
    wire N__5096;
    wire N__5095;
    wire N__5094;
    wire N__5087;
    wire N__5086;
    wire N__5085;
    wire N__5078;
    wire N__5077;
    wire N__5076;
    wire N__5059;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5044;
    wire N__5041;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5029;
    wire N__5026;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5011;
    wire N__5008;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4978;
    wire N__4977;
    wire N__4976;
    wire N__4975;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4953;
    wire N__4952;
    wire N__4951;
    wire N__4950;
    wire N__4949;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4943;
    wire N__4942;
    wire N__4941;
    wire N__4940;
    wire N__4939;
    wire N__4938;
    wire N__4937;
    wire N__4936;
    wire N__4935;
    wire N__4934;
    wire N__4933;
    wire N__4932;
    wire N__4931;
    wire N__4928;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4907;
    wire N__4900;
    wire N__4893;
    wire N__4882;
    wire N__4881;
    wire N__4878;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4862;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4837;
    wire N__4834;
    wire N__4829;
    wire N__4820;
    wire N__4815;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4765;
    wire N__4764;
    wire N__4763;
    wire N__4762;
    wire N__4761;
    wire N__4760;
    wire N__4759;
    wire N__4758;
    wire N__4757;
    wire N__4756;
    wire N__4755;
    wire N__4754;
    wire N__4753;
    wire N__4752;
    wire N__4751;
    wire N__4750;
    wire N__4749;
    wire N__4748;
    wire N__4747;
    wire N__4746;
    wire N__4745;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4695;
    wire N__4694;
    wire N__4693;
    wire N__4692;
    wire N__4689;
    wire N__4688;
    wire N__4685;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4662;
    wire N__4661;
    wire N__4660;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4641;
    wire N__4638;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4614;
    wire N__4609;
    wire N__4606;
    wire N__4601;
    wire N__4598;
    wire N__4593;
    wire N__4588;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4573;
    wire N__4572;
    wire N__4571;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4530;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4524;
    wire N__4517;
    wire N__4512;
    wire N__4511;
    wire N__4510;
    wire N__4509;
    wire N__4508;
    wire N__4503;
    wire N__4500;
    wire N__4499;
    wire N__4498;
    wire N__4497;
    wire N__4494;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4485;
    wire N__4484;
    wire N__4483;
    wire N__4482;
    wire N__4481;
    wire N__4480;
    wire N__4479;
    wire N__4474;
    wire N__4467;
    wire N__4462;
    wire N__4455;
    wire N__4454;
    wire N__4445;
    wire N__4440;
    wire N__4437;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4384;
    wire N__4381;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4369;
    wire N__4366;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4351;
    wire N__4348;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4336;
    wire N__4333;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4321;
    wire N__4318;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4306;
    wire N__4303;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4291;
    wire N__4288;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4276;
    wire N__4273;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4245;
    wire N__4240;
    wire N__4237;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4225;
    wire N__4222;
    wire N__4219;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4204;
    wire N__4201;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4189;
    wire N__4186;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4174;
    wire N__4171;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4156;
    wire N__4153;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4141;
    wire N__4138;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4126;
    wire N__4123;
    wire N__4122;
    wire N__4121;
    wire N__4120;
    wire N__4117;
    wire N__4110;
    wire N__4109;
    wire N__4108;
    wire N__4107;
    wire N__4106;
    wire N__4105;
    wire N__4104;
    wire N__4103;
    wire N__4102;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4084;
    wire N__4077;
    wire N__4074;
    wire N__4067;
    wire N__4060;
    wire N__4059;
    wire N__4058;
    wire N__4055;
    wire N__4054;
    wire N__4053;
    wire N__4052;
    wire N__4047;
    wire N__4044;
    wire N__4037;
    wire N__4034;
    wire N__4027;
    wire N__4024;
    wire N__4023;
    wire N__4022;
    wire N__4019;
    wire N__4014;
    wire N__4011;
    wire N__4010;
    wire N__4009;
    wire N__4008;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3992;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3964;
    wire N__3961;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3934;
    wire N__3933;
    wire N__3932;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3920;
    wire N__3913;
    wire N__3912;
    wire N__3907;
    wire N__3904;
    wire N__3903;
    wire N__3902;
    wire N__3897;
    wire N__3894;
    wire N__3889;
    wire N__3888;
    wire N__3885;
    wire N__3884;
    wire N__3881;
    wire N__3880;
    wire N__3877;
    wire N__3870;
    wire N__3865;
    wire N__3862;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3847;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3832;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3817;
    wire N__3814;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3726;
    wire N__3721;
    wire N__3718;
    wire N__3717;
    wire N__3716;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3687;
    wire N__3684;
    wire N__3683;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3643;
    wire N__3640;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3628;
    wire N__3627;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3619;
    wire N__3618;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3600;
    wire N__3599;
    wire N__3598;
    wire N__3597;
    wire N__3596;
    wire N__3595;
    wire N__3594;
    wire N__3589;
    wire N__3584;
    wire N__3581;
    wire N__3576;
    wire N__3573;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3549;
    wire N__3546;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3536;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3516;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3480;
    wire N__3477;
    wire N__3476;
    wire N__3473;
    wire N__3470;
    wire N__3467;
    wire N__3460;
    wire N__3459;
    wire N__3458;
    wire N__3457;
    wire N__3456;
    wire N__3455;
    wire N__3454;
    wire N__3453;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3427;
    wire N__3426;
    wire N__3425;
    wire N__3422;
    wire N__3421;
    wire N__3418;
    wire N__3415;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3397;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3385;
    wire N__3384;
    wire N__3381;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3370;
    wire N__3369;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3337;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3325;
    wire N__3324;
    wire N__3321;
    wire N__3320;
    wire N__3319;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3289;
    wire N__3288;
    wire N__3287;
    wire N__3286;
    wire N__3285;
    wire N__3284;
    wire N__3283;
    wire N__3276;
    wire N__3267;
    wire N__3262;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3250;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3222;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3198;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3181;
    wire N__3180;
    wire N__3177;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3129;
    wire N__3128;
    wire N__3125;
    wire N__3120;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3099;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3075;
    wire N__3074;
    wire N__3071;
    wire N__3066;
    wire N__3061;
    wire N__3060;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3040;
    wire N__3039;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3012;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2976;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2961;
    wire N__2956;
    wire N__2955;
    wire N__2954;
    wire N__2951;
    wire N__2946;
    wire N__2941;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2933;
    wire N__2932;
    wire N__2927;
    wire N__2922;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2910;
    wire N__2909;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2841;
    wire N__2838;
    wire N__2835;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2785;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2773;
    wire N__2772;
    wire N__2771;
    wire N__2770;
    wire N__2769;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2730;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2698;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2665;
    wire N__2662;
    wire N__2659;
    wire N__2658;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2643;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2616;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2572;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2562;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2545;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2533;
    wire N__2530;
    wire N__2529;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2505;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2490;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2478;
    wire N__2477;
    wire N__2474;
    wire N__2469;
    wire N__2464;
    wire N__2461;
    wire N__2458;
    wire N__2455;
    wire N__2454;
    wire N__2451;
    wire N__2450;
    wire N__2447;
    wire N__2444;
    wire N__2439;
    wire N__2434;
    wire N__2433;
    wire N__2430;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2413;
    wire N__2410;
    wire N__2407;
    wire N__2404;
    wire N__2401;
    wire N__2398;
    wire N__2397;
    wire N__2396;
    wire N__2393;
    wire N__2388;
    wire N__2383;
    wire N__2380;
    wire N__2377;
    wire N__2374;
    wire N__2373;
    wire N__2372;
    wire N__2369;
    wire N__2364;
    wire N__2359;
    wire N__2358;
    wire N__2357;
    wire N__2356;
    wire N__2355;
    wire N__2354;
    wire N__2353;
    wire N__2352;
    wire N__2351;
    wire N__2350;
    wire N__2349;
    wire N__2348;
    wire N__2347;
    wire N__2346;
    wire N__2345;
    wire N__2344;
    wire N__2341;
    wire N__2338;
    wire N__2335;
    wire N__2332;
    wire N__2329;
    wire N__2326;
    wire N__2323;
    wire N__2320;
    wire N__2317;
    wire N__2314;
    wire N__2311;
    wire N__2308;
    wire N__2305;
    wire N__2302;
    wire N__2299;
    wire N__2296;
    wire N__2295;
    wire N__2294;
    wire N__2293;
    wire N__2292;
    wire N__2291;
    wire N__2290;
    wire N__2289;
    wire N__2280;
    wire N__2271;
    wire N__2262;
    wire N__2253;
    wire N__2250;
    wire N__2247;
    wire N__2244;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2227;
    wire N__2222;
    wire N__2215;
    wire N__2206;
    wire N__2197;
    wire N__2194;
    wire N__2191;
    wire N__2188;
    wire N__2185;
    wire N__2182;
    wire N__2179;
    wire N__2178;
    wire N__2175;
    wire N__2172;
    wire N__2167;
    wire N__2164;
    wire N__2161;
    wire N__2158;
    wire N__2155;
    wire N__2152;
    wire N__2149;
    wire N__2146;
    wire N__2143;
    wire N__2140;
    wire N__2137;
    wire N__2134;
    wire N__2131;
    wire N__2128;
    wire N__2125;
    wire N__2122;
    wire N__2119;
    wire N__2116;
    wire N__2113;
    wire N__2110;
    wire N__2107;
    wire N__2104;
    wire N__2101;
    wire N__2100;
    wire N__2099;
    wire N__2098;
    wire N__2089;
    wire N__2086;
    wire N__2083;
    wire N__2080;
    wire N__2077;
    wire N__2074;
    wire N__2071;
    wire N__2068;
    wire N__2065;
    wire VCCG0;
    wire GNDG0;
    wire \reset_cond.M_stage_qZ0Z_1 ;
    wire \reset_cond.M_stage_qZ0Z_0 ;
    wire rst_n_c;
    wire \reset_cond.M_stage_qZ0Z_2 ;
    wire bfn_26_18_0_;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1 ;
    wire bfn_26_19_0_;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1 ;
    wire bfn_26_20_0_;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1 ;
    wire CONSTANT_ONE_NET;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1 ;
    wire bfn_26_21_0_;
    wire un1_M_count_q_axbxc7_m4_0_a2_2_cascade_;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_0 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_2 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_3 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_10 ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_9 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_8 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_4 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_5 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_CO ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_11 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_CO ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_CO ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_CO ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_CO ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_6 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_CO ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_CO ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_7 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_CO ;
    wire sr_chain_latch_e1_i;
    wire un1_M_count_q_axbxc7_m4_0_a2_3;
    wire M_count_qZ0Z_7;
    wire sr_chain_is_sending_0_clk_cascade_;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_1 ;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_2 ;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_3 ;
    wire sr_data_to_send_4;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_4 ;
    wire sr_data_to_send_5;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_5 ;
    wire sr_data_to_send_6;
    wire sr_data_to_send_7;
    wire M_count_qZ0Z_0;
    wire un1_M_count_q_c2_cascade_;
    wire un1_M_count_q_c5_cascade_;
    wire M_count_qZ0Z_6;
    wire un1_M_count_q_c2;
    wire M_count_qZ0Z_4;
    wire un1_M_count_q_c5;
    wire M_count_qZ0Z_5;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_0_and ;
    wire bfn_28_17_0_;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_1_and ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_0 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_2_and ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_1 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_2 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_3 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_4 ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_24 ;
    wire \sr_chain.M_sr_rest_cycles_q_i_24 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_5 ;
    wire sr_chain_un1_M_sr_rest_cycles_q_1_6;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_12 ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_13 ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_14 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_3_and ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_15 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_17 ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_16 ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_18 ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_19 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_4_and ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_23 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_5_and ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_1_6_i ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_22 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_20 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_CO ;
    wire \sr_chain.M_sr_rest_cycles_qZ0Z_21 ;
    wire N_108_g;
    wire M_count_qZ0Z_1;
    wire sr_data_to_send_1;
    wire M_count_qZ0Z_2;
    wire sr_data_to_send_2;
    wire M_count_qZ0Z_3;
    wire sr_chain_is_sending_0_clk;
    wire sr_data_to_send_3;
    wire \sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_ ;
    wire \sr_chain.M_sr_clock_count_qZ1Z_1 ;
    wire \sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_ ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_5_0_0 ;
    wire sr_data_to_send_0;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_0 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_5_0 ;
    wire \sr_chain.M_main_clock_count_d_0_sqmuxa ;
    wire \sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_ ;
    wire \sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401 ;
    wire \sr_chain.M_main_clock_count_d8_0_and ;
    wire bfn_29_18_0_;
    wire \sr_chain.M_main_clock_count_d8_1_and ;
    wire \sr_chain.M_main_clock_count_d8_0 ;
    wire \sr_chain.M_main_clock_count_d8_2_and ;
    wire \sr_chain.M_main_clock_count_d8_1 ;
    wire \sr_chain.M_main_clock_count_d8_3_and ;
    wire \sr_chain.M_main_clock_count_d8_2 ;
    wire \sr_chain.M_main_clock_count_d8_4_and ;
    wire \sr_chain.M_main_clock_count_d8_3 ;
    wire \sr_chain.M_main_clock_count_d8_5_and ;
    wire \sr_chain.M_main_clock_count_d8_4 ;
    wire \sr_chain.M_main_clock_count_q_i_23 ;
    wire \sr_chain.M_main_clock_count_d8_5 ;
    wire \sr_chain.M_main_clock_count_d8 ;
    wire \sr_chain.latch_0_sqmuxa_1 ;
    wire \sr_chain.M_main_clock_count_d8_THRU_CO ;
    wire \sr_chain.M_sr_clock_count_qZ0Z_0 ;
    wire \sr_chain.M_sr_bit_d12_m_0_cascade_ ;
    wire sr_clk_c;
    wire \sr_chain.M_sr_clock_count_qZ0Z_4 ;
    wire \sr_chain.M_sr_clock_count_qZ0Z_2 ;
    wire \sr_chain.un1_M_sr_clock_count_q_1_c2 ;
    wire \sr_chain.M_sr_clock_count_qZ0Z_3 ;
    wire \sr_chain.M_sr_is_sending_q_RNIMJKTZ0 ;
    wire \sr_chain.un1_M_sr_rest_cycles_q_3_0 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_0 ;
    wire bfn_30_15_0_;
    wire \sr_chain.M_main_clock_count_qZ0Z_1 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_0 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_2 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_1 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_3 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_2 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_4 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_3 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_5 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_4 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_6 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_5 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_7 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_6 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_7 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_8 ;
    wire bfn_30_16_0_;
    wire \sr_chain.M_main_clock_count_qZ0Z_9 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_8 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_10 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_9 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_11 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_10 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_12 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_11 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_13 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_12 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_14 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_13 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_15 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_14 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_15 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_16 ;
    wire bfn_30_17_0_;
    wire \sr_chain.M_main_clock_count_qZ0Z_17 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_16 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_18 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_17 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_19 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_18 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_20 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_19 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_21 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_20 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_22 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_21 ;
    wire \sr_chain.M_main_clock_count_qZ0Z_23 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_22 ;
    wire \sr_chain.un1_M_main_clock_count_q_1_cry_23 ;
    wire bfn_30_18_0_;
    wire \sr_chain.M_main_clock_count_qZ0Z_24 ;
    wire \sr_chain.N_44_g ;
    wire \sr_chain.M_sr_bit_d_2_sqmuxa ;
    wire sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO;
    wire sr_data_c;
    wire clk_c_g;
    wire M_reset_cond_out_0;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_6 ;
    wire \sr_chain.un1_M_sr_clock_count_q ;
    wire \sr_chain.M_sr_data_buffer_qZ0Z_7 ;
    wire sr_chain_latch13;
    wire \sr_chain.M_sr_bit_q_3 ;
    wire _gnd_net_;

    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5114),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__5116),
            .DIN(N__5115),
            .DOUT(N__5114),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__5116),
            .PADOUT(N__5115),
            .PADIN(N__5114),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__5105),
            .DIN(N__5104),
            .DOUT(N__5103),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__5105),
            .PADOUT(N__5104),
            .PADIN(N__5103),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sr_clk_obuf_iopad (
            .OE(N__5096),
            .DIN(N__5095),
            .DOUT(N__5094),
            .PACKAGEPIN(sr_clk));
    defparam sr_clk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sr_clk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sr_clk_obuf_preio (
            .PADOEN(N__5096),
            .PADOUT(N__5095),
            .PADIN(N__5094),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3982),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sr_data_obuf_iopad (
            .OE(N__5087),
            .DIN(N__5086),
            .DOUT(N__5085),
            .PACKAGEPIN(sr_data));
    defparam sr_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sr_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sr_data_obuf_preio (
            .PADOEN(N__5087),
            .PADOUT(N__5086),
            .PADIN(N__5085),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4798),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sr_latch_obuf_iopad (
            .OE(N__5078),
            .DIN(N__5077),
            .DOUT(N__5076),
            .PACKAGEPIN(sr_latch));
    defparam sr_latch_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sr_latch_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sr_latch_obuf_preio (
            .PADOEN(N__5078),
            .PADOUT(N__5077),
            .PADIN(N__5076),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2707),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__1177 (
            .O(N__5059),
            .I(N__5055));
    InMux I__1176 (
            .O(N__5058),
            .I(N__5052));
    LocalMux I__1175 (
            .O(N__5055),
            .I(N__5049));
    LocalMux I__1174 (
            .O(N__5052),
            .I(\sr_chain.M_main_clock_count_qZ0Z_20 ));
    Odrv4 I__1173 (
            .O(N__5049),
            .I(\sr_chain.M_main_clock_count_qZ0Z_20 ));
    InMux I__1172 (
            .O(N__5044),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_19 ));
    InMux I__1171 (
            .O(N__5041),
            .I(N__5037));
    InMux I__1170 (
            .O(N__5040),
            .I(N__5034));
    LocalMux I__1169 (
            .O(N__5037),
            .I(\sr_chain.M_main_clock_count_qZ0Z_21 ));
    LocalMux I__1168 (
            .O(N__5034),
            .I(\sr_chain.M_main_clock_count_qZ0Z_21 ));
    InMux I__1167 (
            .O(N__5029),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_20 ));
    CascadeMux I__1166 (
            .O(N__5026),
            .I(N__5022));
    InMux I__1165 (
            .O(N__5025),
            .I(N__5019));
    InMux I__1164 (
            .O(N__5022),
            .I(N__5016));
    LocalMux I__1163 (
            .O(N__5019),
            .I(\sr_chain.M_main_clock_count_qZ0Z_22 ));
    LocalMux I__1162 (
            .O(N__5016),
            .I(\sr_chain.M_main_clock_count_qZ0Z_22 ));
    InMux I__1161 (
            .O(N__5011),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_21 ));
    InMux I__1160 (
            .O(N__5008),
            .I(N__5004));
    InMux I__1159 (
            .O(N__5007),
            .I(N__5001));
    LocalMux I__1158 (
            .O(N__5004),
            .I(\sr_chain.M_main_clock_count_qZ0Z_23 ));
    LocalMux I__1157 (
            .O(N__5001),
            .I(\sr_chain.M_main_clock_count_qZ0Z_23 ));
    InMux I__1156 (
            .O(N__4996),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_22 ));
    InMux I__1155 (
            .O(N__4993),
            .I(bfn_30_18_0_));
    InMux I__1154 (
            .O(N__4990),
            .I(N__4986));
    InMux I__1153 (
            .O(N__4989),
            .I(N__4983));
    LocalMux I__1152 (
            .O(N__4986),
            .I(\sr_chain.M_main_clock_count_qZ0Z_24 ));
    LocalMux I__1151 (
            .O(N__4983),
            .I(\sr_chain.M_main_clock_count_qZ0Z_24 ));
    SRMux I__1150 (
            .O(N__4978),
            .I(N__4966));
    SRMux I__1149 (
            .O(N__4977),
            .I(N__4966));
    SRMux I__1148 (
            .O(N__4976),
            .I(N__4966));
    SRMux I__1147 (
            .O(N__4975),
            .I(N__4966));
    GlobalMux I__1146 (
            .O(N__4966),
            .I(N__4963));
    gio2CtrlBuf I__1145 (
            .O(N__4963),
            .I(\sr_chain.N_44_g ));
    InMux I__1144 (
            .O(N__4960),
            .I(N__4957));
    LocalMux I__1143 (
            .O(N__4957),
            .I(\sr_chain.M_sr_bit_d_2_sqmuxa ));
    InMux I__1142 (
            .O(N__4954),
            .I(N__4946));
    InMux I__1141 (
            .O(N__4953),
            .I(N__4928));
    InMux I__1140 (
            .O(N__4952),
            .I(N__4923));
    InMux I__1139 (
            .O(N__4951),
            .I(N__4923));
    InMux I__1138 (
            .O(N__4950),
            .I(N__4920));
    InMux I__1137 (
            .O(N__4949),
            .I(N__4917));
    LocalMux I__1136 (
            .O(N__4946),
            .I(N__4911));
    InMux I__1135 (
            .O(N__4945),
            .I(N__4908));
    InMux I__1134 (
            .O(N__4944),
            .I(N__4900));
    InMux I__1133 (
            .O(N__4943),
            .I(N__4900));
    InMux I__1132 (
            .O(N__4942),
            .I(N__4900));
    InMux I__1131 (
            .O(N__4941),
            .I(N__4893));
    InMux I__1130 (
            .O(N__4940),
            .I(N__4893));
    InMux I__1129 (
            .O(N__4939),
            .I(N__4893));
    InMux I__1128 (
            .O(N__4938),
            .I(N__4882));
    InMux I__1127 (
            .O(N__4937),
            .I(N__4882));
    InMux I__1126 (
            .O(N__4936),
            .I(N__4882));
    InMux I__1125 (
            .O(N__4935),
            .I(N__4882));
    InMux I__1124 (
            .O(N__4934),
            .I(N__4882));
    InMux I__1123 (
            .O(N__4933),
            .I(N__4878));
    InMux I__1122 (
            .O(N__4932),
            .I(N__4873));
    InMux I__1121 (
            .O(N__4931),
            .I(N__4873));
    LocalMux I__1120 (
            .O(N__4928),
            .I(N__4870));
    LocalMux I__1119 (
            .O(N__4923),
            .I(N__4867));
    LocalMux I__1118 (
            .O(N__4920),
            .I(N__4862));
    LocalMux I__1117 (
            .O(N__4917),
            .I(N__4862));
    InMux I__1116 (
            .O(N__4916),
            .I(N__4855));
    InMux I__1115 (
            .O(N__4915),
            .I(N__4855));
    InMux I__1114 (
            .O(N__4914),
            .I(N__4855));
    Span4Mux_v I__1113 (
            .O(N__4911),
            .I(N__4850));
    LocalMux I__1112 (
            .O(N__4908),
            .I(N__4847));
    InMux I__1111 (
            .O(N__4907),
            .I(N__4844));
    LocalMux I__1110 (
            .O(N__4900),
            .I(N__4837));
    LocalMux I__1109 (
            .O(N__4893),
            .I(N__4837));
    LocalMux I__1108 (
            .O(N__4882),
            .I(N__4837));
    InMux I__1107 (
            .O(N__4881),
            .I(N__4834));
    LocalMux I__1106 (
            .O(N__4878),
            .I(N__4829));
    LocalMux I__1105 (
            .O(N__4873),
            .I(N__4829));
    Span4Mux_v I__1104 (
            .O(N__4870),
            .I(N__4820));
    Span4Mux_v I__1103 (
            .O(N__4867),
            .I(N__4820));
    Span4Mux_v I__1102 (
            .O(N__4862),
            .I(N__4820));
    LocalMux I__1101 (
            .O(N__4855),
            .I(N__4820));
    InMux I__1100 (
            .O(N__4854),
            .I(N__4815));
    InMux I__1099 (
            .O(N__4853),
            .I(N__4815));
    Odrv4 I__1098 (
            .O(N__4850),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    Odrv4 I__1097 (
            .O(N__4847),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    LocalMux I__1096 (
            .O(N__4844),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    Odrv4 I__1095 (
            .O(N__4837),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    LocalMux I__1094 (
            .O(N__4834),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    Odrv12 I__1093 (
            .O(N__4829),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    Odrv4 I__1092 (
            .O(N__4820),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    LocalMux I__1091 (
            .O(N__4815),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO));
    IoInMux I__1090 (
            .O(N__4798),
            .I(N__4795));
    LocalMux I__1089 (
            .O(N__4795),
            .I(N__4792));
    IoSpan4Mux I__1088 (
            .O(N__4792),
            .I(N__4789));
    Span4Mux_s2_h I__1087 (
            .O(N__4789),
            .I(N__4786));
    Sp12to4 I__1086 (
            .O(N__4786),
            .I(N__4783));
    Span12Mux_s10_h I__1085 (
            .O(N__4783),
            .I(N__4779));
    CascadeMux I__1084 (
            .O(N__4782),
            .I(N__4776));
    Span12Mux_h I__1083 (
            .O(N__4779),
            .I(N__4773));
    InMux I__1082 (
            .O(N__4776),
            .I(N__4770));
    Odrv12 I__1081 (
            .O(N__4773),
            .I(sr_data_c));
    LocalMux I__1080 (
            .O(N__4770),
            .I(sr_data_c));
    ClkMux I__1079 (
            .O(N__4765),
            .I(N__4702));
    ClkMux I__1078 (
            .O(N__4764),
            .I(N__4702));
    ClkMux I__1077 (
            .O(N__4763),
            .I(N__4702));
    ClkMux I__1076 (
            .O(N__4762),
            .I(N__4702));
    ClkMux I__1075 (
            .O(N__4761),
            .I(N__4702));
    ClkMux I__1074 (
            .O(N__4760),
            .I(N__4702));
    ClkMux I__1073 (
            .O(N__4759),
            .I(N__4702));
    ClkMux I__1072 (
            .O(N__4758),
            .I(N__4702));
    ClkMux I__1071 (
            .O(N__4757),
            .I(N__4702));
    ClkMux I__1070 (
            .O(N__4756),
            .I(N__4702));
    ClkMux I__1069 (
            .O(N__4755),
            .I(N__4702));
    ClkMux I__1068 (
            .O(N__4754),
            .I(N__4702));
    ClkMux I__1067 (
            .O(N__4753),
            .I(N__4702));
    ClkMux I__1066 (
            .O(N__4752),
            .I(N__4702));
    ClkMux I__1065 (
            .O(N__4751),
            .I(N__4702));
    ClkMux I__1064 (
            .O(N__4750),
            .I(N__4702));
    ClkMux I__1063 (
            .O(N__4749),
            .I(N__4702));
    ClkMux I__1062 (
            .O(N__4748),
            .I(N__4702));
    ClkMux I__1061 (
            .O(N__4747),
            .I(N__4702));
    ClkMux I__1060 (
            .O(N__4746),
            .I(N__4702));
    ClkMux I__1059 (
            .O(N__4745),
            .I(N__4702));
    GlobalMux I__1058 (
            .O(N__4702),
            .I(N__4699));
    gio2CtrlBuf I__1057 (
            .O(N__4699),
            .I(clk_c_g));
    IoInMux I__1056 (
            .O(N__4696),
            .I(N__4689));
    SRMux I__1055 (
            .O(N__4695),
            .I(N__4685));
    SRMux I__1054 (
            .O(N__4694),
            .I(N__4681));
    SRMux I__1053 (
            .O(N__4693),
            .I(N__4678));
    SRMux I__1052 (
            .O(N__4692),
            .I(N__4675));
    LocalMux I__1051 (
            .O(N__4689),
            .I(N__4672));
    SRMux I__1050 (
            .O(N__4688),
            .I(N__4669));
    LocalMux I__1049 (
            .O(N__4685),
            .I(N__4666));
    SRMux I__1048 (
            .O(N__4684),
            .I(N__4663));
    LocalMux I__1047 (
            .O(N__4681),
            .I(N__4655));
    LocalMux I__1046 (
            .O(N__4678),
            .I(N__4655));
    LocalMux I__1045 (
            .O(N__4675),
            .I(N__4652));
    Span4Mux_s1_v I__1044 (
            .O(N__4672),
            .I(N__4649));
    LocalMux I__1043 (
            .O(N__4669),
            .I(N__4646));
    Span4Mux_v I__1042 (
            .O(N__4666),
            .I(N__4641));
    LocalMux I__1041 (
            .O(N__4663),
            .I(N__4641));
    InMux I__1040 (
            .O(N__4662),
            .I(N__4638));
    InMux I__1039 (
            .O(N__4661),
            .I(N__4633));
    InMux I__1038 (
            .O(N__4660),
            .I(N__4633));
    Span4Mux_v I__1037 (
            .O(N__4655),
            .I(N__4630));
    Span4Mux_v I__1036 (
            .O(N__4652),
            .I(N__4627));
    Sp12to4 I__1035 (
            .O(N__4649),
            .I(N__4624));
    Span4Mux_h I__1034 (
            .O(N__4646),
            .I(N__4621));
    Sp12to4 I__1033 (
            .O(N__4641),
            .I(N__4614));
    LocalMux I__1032 (
            .O(N__4638),
            .I(N__4614));
    LocalMux I__1031 (
            .O(N__4633),
            .I(N__4614));
    Span4Mux_h I__1030 (
            .O(N__4630),
            .I(N__4609));
    Span4Mux_h I__1029 (
            .O(N__4627),
            .I(N__4609));
    Span12Mux_h I__1028 (
            .O(N__4624),
            .I(N__4606));
    Sp12to4 I__1027 (
            .O(N__4621),
            .I(N__4601));
    Span12Mux_v I__1026 (
            .O(N__4614),
            .I(N__4601));
    Span4Mux_h I__1025 (
            .O(N__4609),
            .I(N__4598));
    Span12Mux_v I__1024 (
            .O(N__4606),
            .I(N__4593));
    Span12Mux_h I__1023 (
            .O(N__4601),
            .I(N__4593));
    Odrv4 I__1022 (
            .O(N__4598),
            .I(M_reset_cond_out_0));
    Odrv12 I__1021 (
            .O(N__4593),
            .I(M_reset_cond_out_0));
    InMux I__1020 (
            .O(N__4588),
            .I(N__4584));
    InMux I__1019 (
            .O(N__4587),
            .I(N__4581));
    LocalMux I__1018 (
            .O(N__4584),
            .I(N__4578));
    LocalMux I__1017 (
            .O(N__4581),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_6 ));
    Odrv4 I__1016 (
            .O(N__4578),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_6 ));
    CascadeMux I__1015 (
            .O(N__4573),
            .I(N__4567));
    InMux I__1014 (
            .O(N__4572),
            .I(N__4564));
    InMux I__1013 (
            .O(N__4571),
            .I(N__4559));
    InMux I__1012 (
            .O(N__4570),
            .I(N__4559));
    InMux I__1011 (
            .O(N__4567),
            .I(N__4556));
    LocalMux I__1010 (
            .O(N__4564),
            .I(N__4553));
    LocalMux I__1009 (
            .O(N__4559),
            .I(N__4550));
    LocalMux I__1008 (
            .O(N__4556),
            .I(\sr_chain.un1_M_sr_clock_count_q ));
    Odrv4 I__1007 (
            .O(N__4553),
            .I(\sr_chain.un1_M_sr_clock_count_q ));
    Odrv12 I__1006 (
            .O(N__4550),
            .I(\sr_chain.un1_M_sr_clock_count_q ));
    CascadeMux I__1005 (
            .O(N__4543),
            .I(N__4540));
    InMux I__1004 (
            .O(N__4540),
            .I(N__4537));
    LocalMux I__1003 (
            .O(N__4537),
            .I(N__4534));
    Odrv12 I__1002 (
            .O(N__4534),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_7 ));
    CascadeMux I__1001 (
            .O(N__4531),
            .I(N__4525));
    InMux I__1000 (
            .O(N__4530),
            .I(N__4517));
    InMux I__999 (
            .O(N__4529),
            .I(N__4517));
    InMux I__998 (
            .O(N__4528),
            .I(N__4517));
    InMux I__997 (
            .O(N__4525),
            .I(N__4512));
    InMux I__996 (
            .O(N__4524),
            .I(N__4512));
    LocalMux I__995 (
            .O(N__4517),
            .I(N__4503));
    LocalMux I__994 (
            .O(N__4512),
            .I(N__4503));
    InMux I__993 (
            .O(N__4511),
            .I(N__4500));
    CascadeMux I__992 (
            .O(N__4510),
            .I(N__4494));
    CascadeMux I__991 (
            .O(N__4509),
            .I(N__4490));
    CascadeMux I__990 (
            .O(N__4508),
            .I(N__4487));
    Span4Mux_h I__989 (
            .O(N__4503),
            .I(N__4474));
    LocalMux I__988 (
            .O(N__4500),
            .I(N__4474));
    InMux I__987 (
            .O(N__4499),
            .I(N__4467));
    InMux I__986 (
            .O(N__4498),
            .I(N__4467));
    InMux I__985 (
            .O(N__4497),
            .I(N__4467));
    InMux I__984 (
            .O(N__4494),
            .I(N__4462));
    InMux I__983 (
            .O(N__4493),
            .I(N__4462));
    InMux I__982 (
            .O(N__4490),
            .I(N__4455));
    InMux I__981 (
            .O(N__4487),
            .I(N__4455));
    InMux I__980 (
            .O(N__4486),
            .I(N__4455));
    InMux I__979 (
            .O(N__4485),
            .I(N__4445));
    InMux I__978 (
            .O(N__4484),
            .I(N__4445));
    InMux I__977 (
            .O(N__4483),
            .I(N__4445));
    InMux I__976 (
            .O(N__4482),
            .I(N__4445));
    InMux I__975 (
            .O(N__4481),
            .I(N__4440));
    InMux I__974 (
            .O(N__4480),
            .I(N__4440));
    InMux I__973 (
            .O(N__4479),
            .I(N__4437));
    Span4Mux_s3_h I__972 (
            .O(N__4474),
            .I(N__4432));
    LocalMux I__971 (
            .O(N__4467),
            .I(N__4432));
    LocalMux I__970 (
            .O(N__4462),
            .I(N__4429));
    LocalMux I__969 (
            .O(N__4455),
            .I(N__4426));
    InMux I__968 (
            .O(N__4454),
            .I(N__4423));
    LocalMux I__967 (
            .O(N__4445),
            .I(sr_chain_latch13));
    LocalMux I__966 (
            .O(N__4440),
            .I(sr_chain_latch13));
    LocalMux I__965 (
            .O(N__4437),
            .I(sr_chain_latch13));
    Odrv4 I__964 (
            .O(N__4432),
            .I(sr_chain_latch13));
    Odrv4 I__963 (
            .O(N__4429),
            .I(sr_chain_latch13));
    Odrv4 I__962 (
            .O(N__4426),
            .I(sr_chain_latch13));
    LocalMux I__961 (
            .O(N__4423),
            .I(sr_chain_latch13));
    InMux I__960 (
            .O(N__4408),
            .I(N__4405));
    LocalMux I__959 (
            .O(N__4405),
            .I(N__4402));
    Span4Mux_v I__958 (
            .O(N__4402),
            .I(N__4399));
    Odrv4 I__957 (
            .O(N__4399),
            .I(\sr_chain.M_sr_bit_q_3 ));
    InMux I__956 (
            .O(N__4396),
            .I(N__4392));
    InMux I__955 (
            .O(N__4395),
            .I(N__4389));
    LocalMux I__954 (
            .O(N__4392),
            .I(\sr_chain.M_main_clock_count_qZ0Z_12 ));
    LocalMux I__953 (
            .O(N__4389),
            .I(\sr_chain.M_main_clock_count_qZ0Z_12 ));
    InMux I__952 (
            .O(N__4384),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_11 ));
    InMux I__951 (
            .O(N__4381),
            .I(N__4377));
    InMux I__950 (
            .O(N__4380),
            .I(N__4374));
    LocalMux I__949 (
            .O(N__4377),
            .I(\sr_chain.M_main_clock_count_qZ0Z_13 ));
    LocalMux I__948 (
            .O(N__4374),
            .I(\sr_chain.M_main_clock_count_qZ0Z_13 ));
    InMux I__947 (
            .O(N__4369),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_12 ));
    CascadeMux I__946 (
            .O(N__4366),
            .I(N__4362));
    InMux I__945 (
            .O(N__4365),
            .I(N__4359));
    InMux I__944 (
            .O(N__4362),
            .I(N__4356));
    LocalMux I__943 (
            .O(N__4359),
            .I(\sr_chain.M_main_clock_count_qZ0Z_14 ));
    LocalMux I__942 (
            .O(N__4356),
            .I(\sr_chain.M_main_clock_count_qZ0Z_14 ));
    InMux I__941 (
            .O(N__4351),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_13 ));
    InMux I__940 (
            .O(N__4348),
            .I(N__4344));
    InMux I__939 (
            .O(N__4347),
            .I(N__4341));
    LocalMux I__938 (
            .O(N__4344),
            .I(\sr_chain.M_main_clock_count_qZ0Z_15 ));
    LocalMux I__937 (
            .O(N__4341),
            .I(\sr_chain.M_main_clock_count_qZ0Z_15 ));
    InMux I__936 (
            .O(N__4336),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_14 ));
    InMux I__935 (
            .O(N__4333),
            .I(N__4329));
    InMux I__934 (
            .O(N__4332),
            .I(N__4326));
    LocalMux I__933 (
            .O(N__4329),
            .I(\sr_chain.M_main_clock_count_qZ0Z_16 ));
    LocalMux I__932 (
            .O(N__4326),
            .I(\sr_chain.M_main_clock_count_qZ0Z_16 ));
    InMux I__931 (
            .O(N__4321),
            .I(bfn_30_17_0_));
    InMux I__930 (
            .O(N__4318),
            .I(N__4314));
    InMux I__929 (
            .O(N__4317),
            .I(N__4311));
    LocalMux I__928 (
            .O(N__4314),
            .I(\sr_chain.M_main_clock_count_qZ0Z_17 ));
    LocalMux I__927 (
            .O(N__4311),
            .I(\sr_chain.M_main_clock_count_qZ0Z_17 ));
    InMux I__926 (
            .O(N__4306),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_16 ));
    InMux I__925 (
            .O(N__4303),
            .I(N__4299));
    InMux I__924 (
            .O(N__4302),
            .I(N__4296));
    LocalMux I__923 (
            .O(N__4299),
            .I(\sr_chain.M_main_clock_count_qZ0Z_18 ));
    LocalMux I__922 (
            .O(N__4296),
            .I(\sr_chain.M_main_clock_count_qZ0Z_18 ));
    InMux I__921 (
            .O(N__4291),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_17 ));
    InMux I__920 (
            .O(N__4288),
            .I(N__4284));
    InMux I__919 (
            .O(N__4287),
            .I(N__4281));
    LocalMux I__918 (
            .O(N__4284),
            .I(\sr_chain.M_main_clock_count_qZ0Z_19 ));
    LocalMux I__917 (
            .O(N__4281),
            .I(\sr_chain.M_main_clock_count_qZ0Z_19 ));
    InMux I__916 (
            .O(N__4276),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_18 ));
    InMux I__915 (
            .O(N__4273),
            .I(N__4269));
    InMux I__914 (
            .O(N__4272),
            .I(N__4266));
    LocalMux I__913 (
            .O(N__4269),
            .I(\sr_chain.M_main_clock_count_qZ0Z_3 ));
    LocalMux I__912 (
            .O(N__4266),
            .I(\sr_chain.M_main_clock_count_qZ0Z_3 ));
    InMux I__911 (
            .O(N__4261),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_2 ));
    CascadeMux I__910 (
            .O(N__4258),
            .I(N__4255));
    InMux I__909 (
            .O(N__4255),
            .I(N__4251));
    InMux I__908 (
            .O(N__4254),
            .I(N__4248));
    LocalMux I__907 (
            .O(N__4251),
            .I(N__4245));
    LocalMux I__906 (
            .O(N__4248),
            .I(\sr_chain.M_main_clock_count_qZ0Z_4 ));
    Odrv4 I__905 (
            .O(N__4245),
            .I(\sr_chain.M_main_clock_count_qZ0Z_4 ));
    InMux I__904 (
            .O(N__4240),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_3 ));
    InMux I__903 (
            .O(N__4237),
            .I(N__4233));
    InMux I__902 (
            .O(N__4236),
            .I(N__4230));
    LocalMux I__901 (
            .O(N__4233),
            .I(\sr_chain.M_main_clock_count_qZ0Z_5 ));
    LocalMux I__900 (
            .O(N__4230),
            .I(\sr_chain.M_main_clock_count_qZ0Z_5 ));
    InMux I__899 (
            .O(N__4225),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_4 ));
    CascadeMux I__898 (
            .O(N__4222),
            .I(N__4219));
    InMux I__897 (
            .O(N__4219),
            .I(N__4215));
    InMux I__896 (
            .O(N__4218),
            .I(N__4212));
    LocalMux I__895 (
            .O(N__4215),
            .I(N__4209));
    LocalMux I__894 (
            .O(N__4212),
            .I(\sr_chain.M_main_clock_count_qZ0Z_6 ));
    Odrv4 I__893 (
            .O(N__4209),
            .I(\sr_chain.M_main_clock_count_qZ0Z_6 ));
    InMux I__892 (
            .O(N__4204),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_5 ));
    InMux I__891 (
            .O(N__4201),
            .I(N__4197));
    InMux I__890 (
            .O(N__4200),
            .I(N__4194));
    LocalMux I__889 (
            .O(N__4197),
            .I(\sr_chain.M_main_clock_count_qZ0Z_7 ));
    LocalMux I__888 (
            .O(N__4194),
            .I(\sr_chain.M_main_clock_count_qZ0Z_7 ));
    InMux I__887 (
            .O(N__4189),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_6 ));
    InMux I__886 (
            .O(N__4186),
            .I(N__4182));
    InMux I__885 (
            .O(N__4185),
            .I(N__4179));
    LocalMux I__884 (
            .O(N__4182),
            .I(\sr_chain.M_main_clock_count_qZ0Z_8 ));
    LocalMux I__883 (
            .O(N__4179),
            .I(\sr_chain.M_main_clock_count_qZ0Z_8 ));
    InMux I__882 (
            .O(N__4174),
            .I(bfn_30_16_0_));
    CascadeMux I__881 (
            .O(N__4171),
            .I(N__4167));
    InMux I__880 (
            .O(N__4170),
            .I(N__4164));
    InMux I__879 (
            .O(N__4167),
            .I(N__4161));
    LocalMux I__878 (
            .O(N__4164),
            .I(\sr_chain.M_main_clock_count_qZ0Z_9 ));
    LocalMux I__877 (
            .O(N__4161),
            .I(\sr_chain.M_main_clock_count_qZ0Z_9 ));
    InMux I__876 (
            .O(N__4156),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_8 ));
    InMux I__875 (
            .O(N__4153),
            .I(N__4149));
    InMux I__874 (
            .O(N__4152),
            .I(N__4146));
    LocalMux I__873 (
            .O(N__4149),
            .I(\sr_chain.M_main_clock_count_qZ0Z_10 ));
    LocalMux I__872 (
            .O(N__4146),
            .I(\sr_chain.M_main_clock_count_qZ0Z_10 ));
    InMux I__871 (
            .O(N__4141),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_9 ));
    InMux I__870 (
            .O(N__4138),
            .I(N__4134));
    InMux I__869 (
            .O(N__4137),
            .I(N__4131));
    LocalMux I__868 (
            .O(N__4134),
            .I(\sr_chain.M_main_clock_count_qZ0Z_11 ));
    LocalMux I__867 (
            .O(N__4131),
            .I(\sr_chain.M_main_clock_count_qZ0Z_11 ));
    InMux I__866 (
            .O(N__4126),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_10 ));
    InMux I__865 (
            .O(N__4123),
            .I(N__4117));
    InMux I__864 (
            .O(N__4122),
            .I(N__4110));
    InMux I__863 (
            .O(N__4121),
            .I(N__4110));
    InMux I__862 (
            .O(N__4120),
            .I(N__4110));
    LocalMux I__861 (
            .O(N__4117),
            .I(N__4098));
    LocalMux I__860 (
            .O(N__4110),
            .I(N__4095));
    InMux I__859 (
            .O(N__4109),
            .I(N__4084));
    InMux I__858 (
            .O(N__4108),
            .I(N__4084));
    InMux I__857 (
            .O(N__4107),
            .I(N__4084));
    InMux I__856 (
            .O(N__4106),
            .I(N__4084));
    InMux I__855 (
            .O(N__4105),
            .I(N__4084));
    InMux I__854 (
            .O(N__4104),
            .I(N__4077));
    InMux I__853 (
            .O(N__4103),
            .I(N__4077));
    InMux I__852 (
            .O(N__4102),
            .I(N__4077));
    InMux I__851 (
            .O(N__4101),
            .I(N__4074));
    Span4Mux_v I__850 (
            .O(N__4098),
            .I(N__4067));
    Span4Mux_v I__849 (
            .O(N__4095),
            .I(N__4067));
    LocalMux I__848 (
            .O(N__4084),
            .I(N__4067));
    LocalMux I__847 (
            .O(N__4077),
            .I(\sr_chain.latch_0_sqmuxa_1 ));
    LocalMux I__846 (
            .O(N__4074),
            .I(\sr_chain.latch_0_sqmuxa_1 ));
    Odrv4 I__845 (
            .O(N__4067),
            .I(\sr_chain.latch_0_sqmuxa_1 ));
    InMux I__844 (
            .O(N__4060),
            .I(N__4055));
    InMux I__843 (
            .O(N__4059),
            .I(N__4047));
    InMux I__842 (
            .O(N__4058),
            .I(N__4047));
    LocalMux I__841 (
            .O(N__4055),
            .I(N__4044));
    InMux I__840 (
            .O(N__4054),
            .I(N__4037));
    InMux I__839 (
            .O(N__4053),
            .I(N__4037));
    InMux I__838 (
            .O(N__4052),
            .I(N__4037));
    LocalMux I__837 (
            .O(N__4047),
            .I(N__4034));
    Odrv4 I__836 (
            .O(N__4044),
            .I(\sr_chain.M_main_clock_count_d8_THRU_CO ));
    LocalMux I__835 (
            .O(N__4037),
            .I(\sr_chain.M_main_clock_count_d8_THRU_CO ));
    Odrv4 I__834 (
            .O(N__4034),
            .I(\sr_chain.M_main_clock_count_d8_THRU_CO ));
    CascadeMux I__833 (
            .O(N__4027),
            .I(N__4024));
    InMux I__832 (
            .O(N__4024),
            .I(N__4019));
    InMux I__831 (
            .O(N__4023),
            .I(N__4014));
    InMux I__830 (
            .O(N__4022),
            .I(N__4014));
    LocalMux I__829 (
            .O(N__4019),
            .I(N__4011));
    LocalMux I__828 (
            .O(N__4014),
            .I(N__4004));
    Span4Mux_s3_h I__827 (
            .O(N__4011),
            .I(N__4001));
    InMux I__826 (
            .O(N__4010),
            .I(N__3992));
    InMux I__825 (
            .O(N__4009),
            .I(N__3992));
    InMux I__824 (
            .O(N__4008),
            .I(N__3992));
    InMux I__823 (
            .O(N__4007),
            .I(N__3992));
    Odrv12 I__822 (
            .O(N__4004),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_0 ));
    Odrv4 I__821 (
            .O(N__4001),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_0 ));
    LocalMux I__820 (
            .O(N__3992),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_0 ));
    CascadeMux I__819 (
            .O(N__3985),
            .I(\sr_chain.M_sr_bit_d12_m_0_cascade_ ));
    IoInMux I__818 (
            .O(N__3982),
            .I(N__3979));
    LocalMux I__817 (
            .O(N__3979),
            .I(N__3976));
    Span12Mux_s4_h I__816 (
            .O(N__3976),
            .I(N__3973));
    Span12Mux_h I__815 (
            .O(N__3973),
            .I(N__3970));
    Span12Mux_h I__814 (
            .O(N__3970),
            .I(N__3967));
    Odrv12 I__813 (
            .O(N__3967),
            .I(sr_clk_c));
    CascadeMux I__812 (
            .O(N__3964),
            .I(N__3961));
    InMux I__811 (
            .O(N__3961),
            .I(N__3957));
    CascadeMux I__810 (
            .O(N__3960),
            .I(N__3954));
    LocalMux I__809 (
            .O(N__3957),
            .I(N__3951));
    InMux I__808 (
            .O(N__3954),
            .I(N__3947));
    Span4Mux_v I__807 (
            .O(N__3951),
            .I(N__3944));
    InMux I__806 (
            .O(N__3950),
            .I(N__3941));
    LocalMux I__805 (
            .O(N__3947),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_4 ));
    Odrv4 I__804 (
            .O(N__3944),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_4 ));
    LocalMux I__803 (
            .O(N__3941),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_4 ));
    InMux I__802 (
            .O(N__3934),
            .I(N__3928));
    InMux I__801 (
            .O(N__3933),
            .I(N__3925));
    InMux I__800 (
            .O(N__3932),
            .I(N__3920));
    InMux I__799 (
            .O(N__3931),
            .I(N__3920));
    LocalMux I__798 (
            .O(N__3928),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_2 ));
    LocalMux I__797 (
            .O(N__3925),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_2 ));
    LocalMux I__796 (
            .O(N__3920),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_2 ));
    InMux I__795 (
            .O(N__3913),
            .I(N__3907));
    InMux I__794 (
            .O(N__3912),
            .I(N__3907));
    LocalMux I__793 (
            .O(N__3907),
            .I(\sr_chain.un1_M_sr_clock_count_q_1_c2 ));
    InMux I__792 (
            .O(N__3904),
            .I(N__3897));
    InMux I__791 (
            .O(N__3903),
            .I(N__3897));
    InMux I__790 (
            .O(N__3902),
            .I(N__3894));
    LocalMux I__789 (
            .O(N__3897),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_3 ));
    LocalMux I__788 (
            .O(N__3894),
            .I(\sr_chain.M_sr_clock_count_qZ0Z_3 ));
    SRMux I__787 (
            .O(N__3889),
            .I(N__3885));
    CascadeMux I__786 (
            .O(N__3888),
            .I(N__3881));
    LocalMux I__785 (
            .O(N__3885),
            .I(N__3877));
    InMux I__784 (
            .O(N__3884),
            .I(N__3870));
    InMux I__783 (
            .O(N__3881),
            .I(N__3870));
    InMux I__782 (
            .O(N__3880),
            .I(N__3870));
    Span4Mux_s3_h I__781 (
            .O(N__3877),
            .I(N__3865));
    LocalMux I__780 (
            .O(N__3870),
            .I(N__3865));
    Odrv4 I__779 (
            .O(N__3865),
            .I(\sr_chain.M_sr_is_sending_q_RNIMJKTZ0 ));
    CascadeMux I__778 (
            .O(N__3862),
            .I(N__3858));
    InMux I__777 (
            .O(N__3861),
            .I(N__3855));
    InMux I__776 (
            .O(N__3858),
            .I(N__3852));
    LocalMux I__775 (
            .O(N__3855),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_3_0 ));
    LocalMux I__774 (
            .O(N__3852),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_3_0 ));
    InMux I__773 (
            .O(N__3847),
            .I(N__3843));
    InMux I__772 (
            .O(N__3846),
            .I(N__3840));
    LocalMux I__771 (
            .O(N__3843),
            .I(N__3837));
    LocalMux I__770 (
            .O(N__3840),
            .I(\sr_chain.M_main_clock_count_qZ0Z_0 ));
    Odrv4 I__769 (
            .O(N__3837),
            .I(\sr_chain.M_main_clock_count_qZ0Z_0 ));
    CascadeMux I__768 (
            .O(N__3832),
            .I(N__3828));
    InMux I__767 (
            .O(N__3831),
            .I(N__3825));
    InMux I__766 (
            .O(N__3828),
            .I(N__3822));
    LocalMux I__765 (
            .O(N__3825),
            .I(\sr_chain.M_main_clock_count_qZ0Z_1 ));
    LocalMux I__764 (
            .O(N__3822),
            .I(\sr_chain.M_main_clock_count_qZ0Z_1 ));
    InMux I__763 (
            .O(N__3817),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_0 ));
    InMux I__762 (
            .O(N__3814),
            .I(N__3810));
    InMux I__761 (
            .O(N__3813),
            .I(N__3807));
    LocalMux I__760 (
            .O(N__3810),
            .I(\sr_chain.M_main_clock_count_qZ0Z_2 ));
    LocalMux I__759 (
            .O(N__3807),
            .I(\sr_chain.M_main_clock_count_qZ0Z_2 ));
    InMux I__758 (
            .O(N__3802),
            .I(\sr_chain.un1_M_main_clock_count_q_1_cry_1 ));
    CascadeMux I__757 (
            .O(N__3799),
            .I(N__3796));
    InMux I__756 (
            .O(N__3796),
            .I(N__3793));
    LocalMux I__755 (
            .O(N__3793),
            .I(\sr_chain.M_main_clock_count_d8_0_and ));
    CascadeMux I__754 (
            .O(N__3790),
            .I(N__3787));
    InMux I__753 (
            .O(N__3787),
            .I(N__3784));
    LocalMux I__752 (
            .O(N__3784),
            .I(\sr_chain.M_main_clock_count_d8_1_and ));
    CascadeMux I__751 (
            .O(N__3781),
            .I(N__3778));
    InMux I__750 (
            .O(N__3778),
            .I(N__3775));
    LocalMux I__749 (
            .O(N__3775),
            .I(\sr_chain.M_main_clock_count_d8_2_and ));
    CascadeMux I__748 (
            .O(N__3772),
            .I(N__3769));
    InMux I__747 (
            .O(N__3769),
            .I(N__3766));
    LocalMux I__746 (
            .O(N__3766),
            .I(N__3763));
    Odrv4 I__745 (
            .O(N__3763),
            .I(\sr_chain.M_main_clock_count_d8_3_and ));
    CascadeMux I__744 (
            .O(N__3760),
            .I(N__3757));
    InMux I__743 (
            .O(N__3757),
            .I(N__3754));
    LocalMux I__742 (
            .O(N__3754),
            .I(N__3751));
    Odrv12 I__741 (
            .O(N__3751),
            .I(\sr_chain.M_main_clock_count_d8_4_and ));
    CascadeMux I__740 (
            .O(N__3748),
            .I(N__3745));
    InMux I__739 (
            .O(N__3745),
            .I(N__3742));
    LocalMux I__738 (
            .O(N__3742),
            .I(\sr_chain.M_main_clock_count_d8_5_and ));
    CascadeMux I__737 (
            .O(N__3739),
            .I(N__3736));
    InMux I__736 (
            .O(N__3736),
            .I(N__3733));
    LocalMux I__735 (
            .O(N__3733),
            .I(\sr_chain.M_main_clock_count_q_i_23 ));
    InMux I__734 (
            .O(N__3730),
            .I(\sr_chain.M_main_clock_count_d8 ));
    InMux I__733 (
            .O(N__3727),
            .I(N__3721));
    InMux I__732 (
            .O(N__3726),
            .I(N__3721));
    LocalMux I__731 (
            .O(N__3721),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_5_0 ));
    InMux I__730 (
            .O(N__3718),
            .I(N__3709));
    InMux I__729 (
            .O(N__3717),
            .I(N__3709));
    InMux I__728 (
            .O(N__3716),
            .I(N__3709));
    LocalMux I__727 (
            .O(N__3709),
            .I(N__3706));
    Odrv4 I__726 (
            .O(N__3706),
            .I(\sr_chain.M_main_clock_count_d_0_sqmuxa ));
    CascadeMux I__725 (
            .O(N__3703),
            .I(\sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_ ));
    IoInMux I__724 (
            .O(N__3700),
            .I(N__3697));
    LocalMux I__723 (
            .O(N__3697),
            .I(N__3694));
    Odrv4 I__722 (
            .O(N__3694),
            .I(\sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401 ));
    CascadeMux I__721 (
            .O(N__3691),
            .I(\sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_ ));
    CascadeMux I__720 (
            .O(N__3688),
            .I(N__3684));
    InMux I__719 (
            .O(N__3687),
            .I(N__3676));
    InMux I__718 (
            .O(N__3684),
            .I(N__3676));
    InMux I__717 (
            .O(N__3683),
            .I(N__3676));
    LocalMux I__716 (
            .O(N__3676),
            .I(\sr_chain.M_sr_clock_count_qZ1Z_1 ));
    CascadeMux I__715 (
            .O(N__3673),
            .I(\sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_ ));
    CEMux I__714 (
            .O(N__3670),
            .I(N__3667));
    LocalMux I__713 (
            .O(N__3667),
            .I(N__3664));
    Span4Mux_v I__712 (
            .O(N__3664),
            .I(N__3661));
    Odrv4 I__711 (
            .O(N__3661),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_5_0_0 ));
    InMux I__710 (
            .O(N__3658),
            .I(N__3654));
    InMux I__709 (
            .O(N__3657),
            .I(N__3651));
    LocalMux I__708 (
            .O(N__3654),
            .I(N__3648));
    LocalMux I__707 (
            .O(N__3651),
            .I(sr_data_to_send_0));
    Odrv4 I__706 (
            .O(N__3648),
            .I(sr_data_to_send_0));
    CascadeMux I__705 (
            .O(N__3643),
            .I(N__3640));
    InMux I__704 (
            .O(N__3640),
            .I(N__3636));
    InMux I__703 (
            .O(N__3639),
            .I(N__3633));
    LocalMux I__702 (
            .O(N__3636),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_0 ));
    LocalMux I__701 (
            .O(N__3633),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_0 ));
    InMux I__700 (
            .O(N__3628),
            .I(N__3623));
    CascadeMux I__699 (
            .O(N__3627),
            .I(N__3620));
    CascadeMux I__698 (
            .O(N__3626),
            .I(N__3614));
    LocalMux I__697 (
            .O(N__3623),
            .I(N__3611));
    InMux I__696 (
            .O(N__3620),
            .I(N__3600));
    InMux I__695 (
            .O(N__3619),
            .I(N__3600));
    InMux I__694 (
            .O(N__3618),
            .I(N__3600));
    InMux I__693 (
            .O(N__3617),
            .I(N__3600));
    InMux I__692 (
            .O(N__3614),
            .I(N__3600));
    Span4Mux_h I__691 (
            .O(N__3611),
            .I(N__3589));
    LocalMux I__690 (
            .O(N__3600),
            .I(N__3589));
    InMux I__689 (
            .O(N__3599),
            .I(N__3584));
    InMux I__688 (
            .O(N__3598),
            .I(N__3584));
    InMux I__687 (
            .O(N__3597),
            .I(N__3581));
    InMux I__686 (
            .O(N__3596),
            .I(N__3576));
    InMux I__685 (
            .O(N__3595),
            .I(N__3576));
    InMux I__684 (
            .O(N__3594),
            .I(N__3573));
    Odrv4 I__683 (
            .O(N__3589),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_6_i ));
    LocalMux I__682 (
            .O(N__3584),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_6_i ));
    LocalMux I__681 (
            .O(N__3581),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_6_i ));
    LocalMux I__680 (
            .O(N__3576),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_6_i ));
    LocalMux I__679 (
            .O(N__3573),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_6_i ));
    CascadeMux I__678 (
            .O(N__3562),
            .I(N__3559));
    InMux I__677 (
            .O(N__3559),
            .I(N__3556));
    LocalMux I__676 (
            .O(N__3556),
            .I(N__3553));
    Odrv12 I__675 (
            .O(N__3553),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_CO ));
    InMux I__674 (
            .O(N__3550),
            .I(N__3546));
    InMux I__673 (
            .O(N__3549),
            .I(N__3542));
    LocalMux I__672 (
            .O(N__3546),
            .I(N__3539));
    InMux I__671 (
            .O(N__3545),
            .I(N__3536));
    LocalMux I__670 (
            .O(N__3542),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_22 ));
    Odrv4 I__669 (
            .O(N__3539),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_22 ));
    LocalMux I__668 (
            .O(N__3536),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_22 ));
    CascadeMux I__667 (
            .O(N__3529),
            .I(N__3526));
    InMux I__666 (
            .O(N__3526),
            .I(N__3523));
    LocalMux I__665 (
            .O(N__3523),
            .I(N__3520));
    Odrv4 I__664 (
            .O(N__3520),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_CO ));
    InMux I__663 (
            .O(N__3517),
            .I(N__3512));
    CascadeMux I__662 (
            .O(N__3516),
            .I(N__3509));
    InMux I__661 (
            .O(N__3515),
            .I(N__3506));
    LocalMux I__660 (
            .O(N__3512),
            .I(N__3503));
    InMux I__659 (
            .O(N__3509),
            .I(N__3500));
    LocalMux I__658 (
            .O(N__3506),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_20 ));
    Odrv4 I__657 (
            .O(N__3503),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_20 ));
    LocalMux I__656 (
            .O(N__3500),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_20 ));
    CascadeMux I__655 (
            .O(N__3493),
            .I(N__3490));
    InMux I__654 (
            .O(N__3490),
            .I(N__3487));
    LocalMux I__653 (
            .O(N__3487),
            .I(N__3484));
    Odrv4 I__652 (
            .O(N__3484),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_CO ));
    InMux I__651 (
            .O(N__3481),
            .I(N__3477));
    InMux I__650 (
            .O(N__3480),
            .I(N__3473));
    LocalMux I__649 (
            .O(N__3477),
            .I(N__3470));
    InMux I__648 (
            .O(N__3476),
            .I(N__3467));
    LocalMux I__647 (
            .O(N__3473),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_21 ));
    Odrv4 I__646 (
            .O(N__3470),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_21 ));
    LocalMux I__645 (
            .O(N__3467),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_21 ));
    SRMux I__644 (
            .O(N__3460),
            .I(N__3436));
    SRMux I__643 (
            .O(N__3459),
            .I(N__3436));
    SRMux I__642 (
            .O(N__3458),
            .I(N__3436));
    SRMux I__641 (
            .O(N__3457),
            .I(N__3436));
    SRMux I__640 (
            .O(N__3456),
            .I(N__3436));
    SRMux I__639 (
            .O(N__3455),
            .I(N__3436));
    SRMux I__638 (
            .O(N__3454),
            .I(N__3436));
    SRMux I__637 (
            .O(N__3453),
            .I(N__3436));
    GlobalMux I__636 (
            .O(N__3436),
            .I(N__3433));
    gio2CtrlBuf I__635 (
            .O(N__3433),
            .I(N_108_g));
    InMux I__634 (
            .O(N__3430),
            .I(N__3427));
    LocalMux I__633 (
            .O(N__3427),
            .I(N__3422));
    CascadeMux I__632 (
            .O(N__3426),
            .I(N__3418));
    InMux I__631 (
            .O(N__3425),
            .I(N__3415));
    Span4Mux_v I__630 (
            .O(N__3422),
            .I(N__3412));
    InMux I__629 (
            .O(N__3421),
            .I(N__3409));
    InMux I__628 (
            .O(N__3418),
            .I(N__3406));
    LocalMux I__627 (
            .O(N__3415),
            .I(M_count_qZ0Z_1));
    Odrv4 I__626 (
            .O(N__3412),
            .I(M_count_qZ0Z_1));
    LocalMux I__625 (
            .O(N__3409),
            .I(M_count_qZ0Z_1));
    LocalMux I__624 (
            .O(N__3406),
            .I(M_count_qZ0Z_1));
    InMux I__623 (
            .O(N__3397),
            .I(N__3393));
    InMux I__622 (
            .O(N__3396),
            .I(N__3390));
    LocalMux I__621 (
            .O(N__3393),
            .I(sr_data_to_send_1));
    LocalMux I__620 (
            .O(N__3390),
            .I(sr_data_to_send_1));
    CascadeMux I__619 (
            .O(N__3385),
            .I(N__3381));
    InMux I__618 (
            .O(N__3384),
            .I(N__3377));
    InMux I__617 (
            .O(N__3381),
            .I(N__3374));
    CascadeMux I__616 (
            .O(N__3380),
            .I(N__3371));
    LocalMux I__615 (
            .O(N__3377),
            .I(N__3365));
    LocalMux I__614 (
            .O(N__3374),
            .I(N__3362));
    InMux I__613 (
            .O(N__3371),
            .I(N__3357));
    InMux I__612 (
            .O(N__3370),
            .I(N__3357));
    InMux I__611 (
            .O(N__3369),
            .I(N__3354));
    InMux I__610 (
            .O(N__3368),
            .I(N__3351));
    Span4Mux_h I__609 (
            .O(N__3365),
            .I(N__3348));
    Odrv4 I__608 (
            .O(N__3362),
            .I(M_count_qZ0Z_2));
    LocalMux I__607 (
            .O(N__3357),
            .I(M_count_qZ0Z_2));
    LocalMux I__606 (
            .O(N__3354),
            .I(M_count_qZ0Z_2));
    LocalMux I__605 (
            .O(N__3351),
            .I(M_count_qZ0Z_2));
    Odrv4 I__604 (
            .O(N__3348),
            .I(M_count_qZ0Z_2));
    InMux I__603 (
            .O(N__3337),
            .I(N__3333));
    InMux I__602 (
            .O(N__3336),
            .I(N__3330));
    LocalMux I__601 (
            .O(N__3333),
            .I(sr_data_to_send_2));
    LocalMux I__600 (
            .O(N__3330),
            .I(sr_data_to_send_2));
    InMux I__599 (
            .O(N__3325),
            .I(N__3321));
    CascadeMux I__598 (
            .O(N__3324),
            .I(N__3315));
    LocalMux I__597 (
            .O(N__3321),
            .I(N__3312));
    InMux I__596 (
            .O(N__3320),
            .I(N__3309));
    InMux I__595 (
            .O(N__3319),
            .I(N__3304));
    InMux I__594 (
            .O(N__3318),
            .I(N__3304));
    InMux I__593 (
            .O(N__3315),
            .I(N__3301));
    Span4Mux_h I__592 (
            .O(N__3312),
            .I(N__3298));
    LocalMux I__591 (
            .O(N__3309),
            .I(M_count_qZ0Z_3));
    LocalMux I__590 (
            .O(N__3304),
            .I(M_count_qZ0Z_3));
    LocalMux I__589 (
            .O(N__3301),
            .I(M_count_qZ0Z_3));
    Odrv4 I__588 (
            .O(N__3298),
            .I(M_count_qZ0Z_3));
    InMux I__587 (
            .O(N__3289),
            .I(N__3276));
    InMux I__586 (
            .O(N__3288),
            .I(N__3276));
    InMux I__585 (
            .O(N__3287),
            .I(N__3276));
    InMux I__584 (
            .O(N__3286),
            .I(N__3267));
    InMux I__583 (
            .O(N__3285),
            .I(N__3267));
    InMux I__582 (
            .O(N__3284),
            .I(N__3267));
    InMux I__581 (
            .O(N__3283),
            .I(N__3267));
    LocalMux I__580 (
            .O(N__3276),
            .I(sr_chain_is_sending_0_clk));
    LocalMux I__579 (
            .O(N__3267),
            .I(sr_chain_is_sending_0_clk));
    InMux I__578 (
            .O(N__3262),
            .I(N__3258));
    InMux I__577 (
            .O(N__3261),
            .I(N__3255));
    LocalMux I__576 (
            .O(N__3258),
            .I(sr_data_to_send_3));
    LocalMux I__575 (
            .O(N__3255),
            .I(sr_data_to_send_3));
    InMux I__574 (
            .O(N__3250),
            .I(N__3246));
    InMux I__573 (
            .O(N__3249),
            .I(N__3243));
    LocalMux I__572 (
            .O(N__3246),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_24 ));
    LocalMux I__571 (
            .O(N__3243),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_24 ));
    CascadeMux I__570 (
            .O(N__3238),
            .I(N__3235));
    InMux I__569 (
            .O(N__3235),
            .I(N__3232));
    LocalMux I__568 (
            .O(N__3232),
            .I(\sr_chain.M_sr_rest_cycles_q_i_24 ));
    InMux I__567 (
            .O(N__3229),
            .I(sr_chain_un1_M_sr_rest_cycles_q_1_6));
    CascadeMux I__566 (
            .O(N__3226),
            .I(N__3223));
    InMux I__565 (
            .O(N__3223),
            .I(N__3218));
    InMux I__564 (
            .O(N__3222),
            .I(N__3215));
    InMux I__563 (
            .O(N__3221),
            .I(N__3212));
    LocalMux I__562 (
            .O(N__3218),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_12 ));
    LocalMux I__561 (
            .O(N__3215),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_12 ));
    LocalMux I__560 (
            .O(N__3212),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_12 ));
    CascadeMux I__559 (
            .O(N__3205),
            .I(N__3202));
    InMux I__558 (
            .O(N__3202),
            .I(N__3199));
    LocalMux I__557 (
            .O(N__3199),
            .I(N__3194));
    InMux I__556 (
            .O(N__3198),
            .I(N__3191));
    InMux I__555 (
            .O(N__3197),
            .I(N__3188));
    Odrv4 I__554 (
            .O(N__3194),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_13 ));
    LocalMux I__553 (
            .O(N__3191),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_13 ));
    LocalMux I__552 (
            .O(N__3188),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_13 ));
    CascadeMux I__551 (
            .O(N__3181),
            .I(N__3177));
    CascadeMux I__550 (
            .O(N__3180),
            .I(N__3173));
    InMux I__549 (
            .O(N__3177),
            .I(N__3170));
    InMux I__548 (
            .O(N__3176),
            .I(N__3167));
    InMux I__547 (
            .O(N__3173),
            .I(N__3164));
    LocalMux I__546 (
            .O(N__3170),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_14 ));
    LocalMux I__545 (
            .O(N__3167),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_14 ));
    LocalMux I__544 (
            .O(N__3164),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_14 ));
    CascadeMux I__543 (
            .O(N__3157),
            .I(N__3154));
    InMux I__542 (
            .O(N__3154),
            .I(N__3151));
    LocalMux I__541 (
            .O(N__3151),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_3_and ));
    InMux I__540 (
            .O(N__3148),
            .I(N__3145));
    LocalMux I__539 (
            .O(N__3145),
            .I(N__3142));
    Span4Mux_h I__538 (
            .O(N__3142),
            .I(N__3139));
    Odrv4 I__537 (
            .O(N__3139),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_CO ));
    InMux I__536 (
            .O(N__3136),
            .I(N__3133));
    LocalMux I__535 (
            .O(N__3133),
            .I(N__3130));
    Span4Mux_h I__534 (
            .O(N__3130),
            .I(N__3125));
    InMux I__533 (
            .O(N__3129),
            .I(N__3120));
    InMux I__532 (
            .O(N__3128),
            .I(N__3120));
    Odrv4 I__531 (
            .O(N__3125),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_15 ));
    LocalMux I__530 (
            .O(N__3120),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_15 ));
    CascadeMux I__529 (
            .O(N__3115),
            .I(N__3112));
    InMux I__528 (
            .O(N__3112),
            .I(N__3109));
    LocalMux I__527 (
            .O(N__3109),
            .I(N__3106));
    Span4Mux_h I__526 (
            .O(N__3106),
            .I(N__3103));
    Odrv4 I__525 (
            .O(N__3103),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_CO ));
    InMux I__524 (
            .O(N__3100),
            .I(N__3095));
    InMux I__523 (
            .O(N__3099),
            .I(N__3092));
    InMux I__522 (
            .O(N__3098),
            .I(N__3089));
    LocalMux I__521 (
            .O(N__3095),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_17 ));
    LocalMux I__520 (
            .O(N__3092),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_17 ));
    LocalMux I__519 (
            .O(N__3089),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_17 ));
    InMux I__518 (
            .O(N__3082),
            .I(N__3079));
    LocalMux I__517 (
            .O(N__3079),
            .I(N__3076));
    Span4Mux_h I__516 (
            .O(N__3076),
            .I(N__3071));
    InMux I__515 (
            .O(N__3075),
            .I(N__3066));
    InMux I__514 (
            .O(N__3074),
            .I(N__3066));
    Odrv4 I__513 (
            .O(N__3071),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_16 ));
    LocalMux I__512 (
            .O(N__3066),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_16 ));
    CascadeMux I__511 (
            .O(N__3061),
            .I(N__3056));
    InMux I__510 (
            .O(N__3060),
            .I(N__3053));
    InMux I__509 (
            .O(N__3059),
            .I(N__3050));
    InMux I__508 (
            .O(N__3056),
            .I(N__3047));
    LocalMux I__507 (
            .O(N__3053),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_18 ));
    LocalMux I__506 (
            .O(N__3050),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_18 ));
    LocalMux I__505 (
            .O(N__3047),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_18 ));
    InMux I__504 (
            .O(N__3040),
            .I(N__3035));
    InMux I__503 (
            .O(N__3039),
            .I(N__3032));
    InMux I__502 (
            .O(N__3038),
            .I(N__3029));
    LocalMux I__501 (
            .O(N__3035),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_19 ));
    LocalMux I__500 (
            .O(N__3032),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_19 ));
    LocalMux I__499 (
            .O(N__3029),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_19 ));
    CascadeMux I__498 (
            .O(N__3022),
            .I(N__3019));
    InMux I__497 (
            .O(N__3019),
            .I(N__3016));
    LocalMux I__496 (
            .O(N__3016),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_4_and ));
    InMux I__495 (
            .O(N__3013),
            .I(N__3008));
    InMux I__494 (
            .O(N__3012),
            .I(N__3005));
    InMux I__493 (
            .O(N__3011),
            .I(N__3002));
    LocalMux I__492 (
            .O(N__3008),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_23 ));
    LocalMux I__491 (
            .O(N__3005),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_23 ));
    LocalMux I__490 (
            .O(N__3002),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_23 ));
    CascadeMux I__489 (
            .O(N__2995),
            .I(N__2992));
    InMux I__488 (
            .O(N__2992),
            .I(N__2989));
    LocalMux I__487 (
            .O(N__2989),
            .I(N__2986));
    Odrv4 I__486 (
            .O(N__2986),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_5_and ));
    CascadeMux I__485 (
            .O(N__2983),
            .I(un1_M_count_q_c2_cascade_));
    CascadeMux I__484 (
            .O(N__2980),
            .I(un1_M_count_q_c5_cascade_));
    InMux I__483 (
            .O(N__2977),
            .I(N__2972));
    InMux I__482 (
            .O(N__2976),
            .I(N__2969));
    InMux I__481 (
            .O(N__2975),
            .I(N__2966));
    LocalMux I__480 (
            .O(N__2972),
            .I(N__2961));
    LocalMux I__479 (
            .O(N__2969),
            .I(N__2961));
    LocalMux I__478 (
            .O(N__2966),
            .I(M_count_qZ0Z_6));
    Odrv4 I__477 (
            .O(N__2961),
            .I(M_count_qZ0Z_6));
    InMux I__476 (
            .O(N__2956),
            .I(N__2951));
    InMux I__475 (
            .O(N__2955),
            .I(N__2946));
    InMux I__474 (
            .O(N__2954),
            .I(N__2946));
    LocalMux I__473 (
            .O(N__2951),
            .I(un1_M_count_q_c2));
    LocalMux I__472 (
            .O(N__2946),
            .I(un1_M_count_q_c2));
    InMux I__471 (
            .O(N__2941),
            .I(N__2937));
    InMux I__470 (
            .O(N__2940),
            .I(N__2934));
    LocalMux I__469 (
            .O(N__2937),
            .I(N__2927));
    LocalMux I__468 (
            .O(N__2934),
            .I(N__2927));
    InMux I__467 (
            .O(N__2933),
            .I(N__2922));
    InMux I__466 (
            .O(N__2932),
            .I(N__2922));
    Odrv4 I__465 (
            .O(N__2927),
            .I(M_count_qZ0Z_4));
    LocalMux I__464 (
            .O(N__2922),
            .I(M_count_qZ0Z_4));
    InMux I__463 (
            .O(N__2917),
            .I(N__2914));
    LocalMux I__462 (
            .O(N__2914),
            .I(un1_M_count_q_c5));
    InMux I__461 (
            .O(N__2911),
            .I(N__2905));
    InMux I__460 (
            .O(N__2910),
            .I(N__2902));
    InMux I__459 (
            .O(N__2909),
            .I(N__2897));
    InMux I__458 (
            .O(N__2908),
            .I(N__2897));
    LocalMux I__457 (
            .O(N__2905),
            .I(N__2894));
    LocalMux I__456 (
            .O(N__2902),
            .I(N__2891));
    LocalMux I__455 (
            .O(N__2897),
            .I(M_count_qZ0Z_5));
    Odrv4 I__454 (
            .O(N__2894),
            .I(M_count_qZ0Z_5));
    Odrv4 I__453 (
            .O(N__2891),
            .I(M_count_qZ0Z_5));
    CascadeMux I__452 (
            .O(N__2884),
            .I(N__2881));
    InMux I__451 (
            .O(N__2881),
            .I(N__2878));
    LocalMux I__450 (
            .O(N__2878),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_0_and ));
    InMux I__449 (
            .O(N__2875),
            .I(N__2872));
    LocalMux I__448 (
            .O(N__2872),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_1_and ));
    InMux I__447 (
            .O(N__2869),
            .I(N__2866));
    LocalMux I__446 (
            .O(N__2866),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_1_2_and ));
    CascadeMux I__445 (
            .O(N__2863),
            .I(sr_chain_is_sending_0_clk_cascade_));
    InMux I__444 (
            .O(N__2860),
            .I(N__2857));
    LocalMux I__443 (
            .O(N__2857),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_1 ));
    InMux I__442 (
            .O(N__2854),
            .I(N__2851));
    LocalMux I__441 (
            .O(N__2851),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_2 ));
    InMux I__440 (
            .O(N__2848),
            .I(N__2845));
    LocalMux I__439 (
            .O(N__2845),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_3 ));
    InMux I__438 (
            .O(N__2842),
            .I(N__2838));
    InMux I__437 (
            .O(N__2841),
            .I(N__2835));
    LocalMux I__436 (
            .O(N__2838),
            .I(sr_data_to_send_4));
    LocalMux I__435 (
            .O(N__2835),
            .I(sr_data_to_send_4));
    InMux I__434 (
            .O(N__2830),
            .I(N__2827));
    LocalMux I__433 (
            .O(N__2827),
            .I(N__2824));
    Odrv4 I__432 (
            .O(N__2824),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_4 ));
    CascadeMux I__431 (
            .O(N__2821),
            .I(N__2818));
    InMux I__430 (
            .O(N__2818),
            .I(N__2814));
    InMux I__429 (
            .O(N__2817),
            .I(N__2811));
    LocalMux I__428 (
            .O(N__2814),
            .I(sr_data_to_send_5));
    LocalMux I__427 (
            .O(N__2811),
            .I(sr_data_to_send_5));
    InMux I__426 (
            .O(N__2806),
            .I(N__2803));
    LocalMux I__425 (
            .O(N__2803),
            .I(N__2800));
    Odrv4 I__424 (
            .O(N__2800),
            .I(\sr_chain.M_sr_data_buffer_qZ0Z_5 ));
    InMux I__423 (
            .O(N__2797),
            .I(N__2793));
    InMux I__422 (
            .O(N__2796),
            .I(N__2790));
    LocalMux I__421 (
            .O(N__2793),
            .I(sr_data_to_send_6));
    LocalMux I__420 (
            .O(N__2790),
            .I(sr_data_to_send_6));
    InMux I__419 (
            .O(N__2785),
            .I(N__2781));
    InMux I__418 (
            .O(N__2784),
            .I(N__2778));
    LocalMux I__417 (
            .O(N__2781),
            .I(sr_data_to_send_7));
    LocalMux I__416 (
            .O(N__2778),
            .I(sr_data_to_send_7));
    InMux I__415 (
            .O(N__2773),
            .I(N__2764));
    InMux I__414 (
            .O(N__2772),
            .I(N__2764));
    InMux I__413 (
            .O(N__2771),
            .I(N__2761));
    InMux I__412 (
            .O(N__2770),
            .I(N__2758));
    InMux I__411 (
            .O(N__2769),
            .I(N__2755));
    LocalMux I__410 (
            .O(N__2764),
            .I(M_count_qZ0Z_0));
    LocalMux I__409 (
            .O(N__2761),
            .I(M_count_qZ0Z_0));
    LocalMux I__408 (
            .O(N__2758),
            .I(M_count_qZ0Z_0));
    LocalMux I__407 (
            .O(N__2755),
            .I(M_count_qZ0Z_0));
    CascadeMux I__406 (
            .O(N__2746),
            .I(N__2743));
    InMux I__405 (
            .O(N__2743),
            .I(N__2740));
    LocalMux I__404 (
            .O(N__2740),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_CO ));
    InMux I__403 (
            .O(N__2737),
            .I(N__2734));
    LocalMux I__402 (
            .O(N__2734),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_CO ));
    InMux I__401 (
            .O(N__2731),
            .I(N__2726));
    InMux I__400 (
            .O(N__2730),
            .I(N__2723));
    InMux I__399 (
            .O(N__2729),
            .I(N__2720));
    LocalMux I__398 (
            .O(N__2726),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_7 ));
    LocalMux I__397 (
            .O(N__2723),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_7 ));
    LocalMux I__396 (
            .O(N__2720),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_7 ));
    InMux I__395 (
            .O(N__2713),
            .I(N__2710));
    LocalMux I__394 (
            .O(N__2710),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_CO ));
    IoInMux I__393 (
            .O(N__2707),
            .I(N__2704));
    LocalMux I__392 (
            .O(N__2704),
            .I(N__2701));
    Span4Mux_s1_h I__391 (
            .O(N__2701),
            .I(N__2698));
    Sp12to4 I__390 (
            .O(N__2698),
            .I(N__2695));
    Span12Mux_s11_v I__389 (
            .O(N__2695),
            .I(N__2692));
    Span12Mux_h I__388 (
            .O(N__2692),
            .I(N__2689));
    Span12Mux_h I__387 (
            .O(N__2689),
            .I(N__2686));
    Odrv12 I__386 (
            .O(N__2686),
            .I(sr_chain_latch_e1_i));
    InMux I__385 (
            .O(N__2683),
            .I(N__2680));
    LocalMux I__384 (
            .O(N__2680),
            .I(un1_M_count_q_axbxc7_m4_0_a2_3));
    InMux I__383 (
            .O(N__2677),
            .I(N__2673));
    InMux I__382 (
            .O(N__2676),
            .I(N__2670));
    LocalMux I__381 (
            .O(N__2673),
            .I(M_count_qZ0Z_7));
    LocalMux I__380 (
            .O(N__2670),
            .I(M_count_qZ0Z_7));
    InMux I__379 (
            .O(N__2665),
            .I(N__2662));
    LocalMux I__378 (
            .O(N__2662),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_CO ));
    CascadeMux I__377 (
            .O(N__2659),
            .I(N__2654));
    CascadeMux I__376 (
            .O(N__2658),
            .I(N__2651));
    InMux I__375 (
            .O(N__2657),
            .I(N__2648));
    InMux I__374 (
            .O(N__2654),
            .I(N__2643));
    InMux I__373 (
            .O(N__2651),
            .I(N__2643));
    LocalMux I__372 (
            .O(N__2648),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_5 ));
    LocalMux I__371 (
            .O(N__2643),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_5 ));
    CascadeMux I__370 (
            .O(N__2638),
            .I(N__2635));
    InMux I__369 (
            .O(N__2635),
            .I(N__2632));
    LocalMux I__368 (
            .O(N__2632),
            .I(N__2629));
    Odrv4 I__367 (
            .O(N__2629),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_CO ));
    CascadeMux I__366 (
            .O(N__2626),
            .I(N__2623));
    InMux I__365 (
            .O(N__2623),
            .I(N__2620));
    LocalMux I__364 (
            .O(N__2620),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_CO ));
    InMux I__363 (
            .O(N__2617),
            .I(N__2612));
    InMux I__362 (
            .O(N__2616),
            .I(N__2609));
    InMux I__361 (
            .O(N__2615),
            .I(N__2606));
    LocalMux I__360 (
            .O(N__2612),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_11 ));
    LocalMux I__359 (
            .O(N__2609),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_11 ));
    LocalMux I__358 (
            .O(N__2606),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_11 ));
    InMux I__357 (
            .O(N__2599),
            .I(N__2596));
    LocalMux I__356 (
            .O(N__2596),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_CO ));
    InMux I__355 (
            .O(N__2593),
            .I(N__2590));
    LocalMux I__354 (
            .O(N__2590),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_CO ));
    InMux I__353 (
            .O(N__2587),
            .I(N__2584));
    LocalMux I__352 (
            .O(N__2584),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_CO ));
    InMux I__351 (
            .O(N__2581),
            .I(N__2578));
    LocalMux I__350 (
            .O(N__2578),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_CO ));
    CascadeMux I__349 (
            .O(N__2575),
            .I(N__2572));
    InMux I__348 (
            .O(N__2572),
            .I(N__2569));
    LocalMux I__347 (
            .O(N__2569),
            .I(N__2566));
    Odrv4 I__346 (
            .O(N__2566),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_CO ));
    InMux I__345 (
            .O(N__2563),
            .I(N__2558));
    InMux I__344 (
            .O(N__2562),
            .I(N__2555));
    InMux I__343 (
            .O(N__2561),
            .I(N__2552));
    LocalMux I__342 (
            .O(N__2558),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_6 ));
    LocalMux I__341 (
            .O(N__2555),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_6 ));
    LocalMux I__340 (
            .O(N__2552),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_6 ));
    CascadeMux I__339 (
            .O(N__2545),
            .I(N__2542));
    InMux I__338 (
            .O(N__2542),
            .I(N__2539));
    LocalMux I__337 (
            .O(N__2539),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_CO ));
    InMux I__336 (
            .O(N__2536),
            .I(N__2533));
    LocalMux I__335 (
            .O(N__2533),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_CO ));
    InMux I__334 (
            .O(N__2530),
            .I(N__2525));
    InMux I__333 (
            .O(N__2529),
            .I(N__2522));
    InMux I__332 (
            .O(N__2528),
            .I(N__2519));
    LocalMux I__331 (
            .O(N__2525),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_1 ));
    LocalMux I__330 (
            .O(N__2522),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_1 ));
    LocalMux I__329 (
            .O(N__2519),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_1 ));
    InMux I__328 (
            .O(N__2512),
            .I(N__2509));
    LocalMux I__327 (
            .O(N__2509),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_CO ));
    CascadeMux I__326 (
            .O(N__2506),
            .I(N__2501));
    CascadeMux I__325 (
            .O(N__2505),
            .I(N__2498));
    InMux I__324 (
            .O(N__2504),
            .I(N__2495));
    InMux I__323 (
            .O(N__2501),
            .I(N__2490));
    InMux I__322 (
            .O(N__2498),
            .I(N__2490));
    LocalMux I__321 (
            .O(N__2495),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_2 ));
    LocalMux I__320 (
            .O(N__2490),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_2 ));
    InMux I__319 (
            .O(N__2485),
            .I(N__2482));
    LocalMux I__318 (
            .O(N__2482),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_CO ));
    InMux I__317 (
            .O(N__2479),
            .I(N__2474));
    InMux I__316 (
            .O(N__2478),
            .I(N__2469));
    InMux I__315 (
            .O(N__2477),
            .I(N__2469));
    LocalMux I__314 (
            .O(N__2474),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_3 ));
    LocalMux I__313 (
            .O(N__2469),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_3 ));
    InMux I__312 (
            .O(N__2464),
            .I(N__2461));
    LocalMux I__311 (
            .O(N__2461),
            .I(N__2458));
    Odrv4 I__310 (
            .O(N__2458),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_CO ));
    InMux I__309 (
            .O(N__2455),
            .I(N__2451));
    CascadeMux I__308 (
            .O(N__2454),
            .I(N__2447));
    LocalMux I__307 (
            .O(N__2451),
            .I(N__2444));
    InMux I__306 (
            .O(N__2450),
            .I(N__2439));
    InMux I__305 (
            .O(N__2447),
            .I(N__2439));
    Odrv4 I__304 (
            .O(N__2444),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_10 ));
    LocalMux I__303 (
            .O(N__2439),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_10 ));
    InMux I__302 (
            .O(N__2434),
            .I(N__2430));
    InMux I__301 (
            .O(N__2433),
            .I(N__2426));
    LocalMux I__300 (
            .O(N__2430),
            .I(N__2423));
    InMux I__299 (
            .O(N__2429),
            .I(N__2420));
    LocalMux I__298 (
            .O(N__2426),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_9 ));
    Odrv4 I__297 (
            .O(N__2423),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_9 ));
    LocalMux I__296 (
            .O(N__2420),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_9 ));
    InMux I__295 (
            .O(N__2413),
            .I(N__2410));
    LocalMux I__294 (
            .O(N__2410),
            .I(N__2407));
    Span4Mux_h I__293 (
            .O(N__2407),
            .I(N__2404));
    Odrv4 I__292 (
            .O(N__2404),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_CO ));
    InMux I__291 (
            .O(N__2401),
            .I(N__2398));
    LocalMux I__290 (
            .O(N__2398),
            .I(N__2393));
    InMux I__289 (
            .O(N__2397),
            .I(N__2388));
    InMux I__288 (
            .O(N__2396),
            .I(N__2388));
    Odrv4 I__287 (
            .O(N__2393),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_8 ));
    LocalMux I__286 (
            .O(N__2388),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_8 ));
    CascadeMux I__285 (
            .O(N__2383),
            .I(N__2380));
    InMux I__284 (
            .O(N__2380),
            .I(N__2377));
    LocalMux I__283 (
            .O(N__2377),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_CO ));
    InMux I__282 (
            .O(N__2374),
            .I(N__2369));
    InMux I__281 (
            .O(N__2373),
            .I(N__2364));
    InMux I__280 (
            .O(N__2372),
            .I(N__2364));
    LocalMux I__279 (
            .O(N__2369),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_4 ));
    LocalMux I__278 (
            .O(N__2364),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_4 ));
    CascadeMux I__277 (
            .O(N__2359),
            .I(N__2341));
    CascadeMux I__276 (
            .O(N__2358),
            .I(N__2338));
    CascadeMux I__275 (
            .O(N__2357),
            .I(N__2335));
    CascadeMux I__274 (
            .O(N__2356),
            .I(N__2332));
    CascadeMux I__273 (
            .O(N__2355),
            .I(N__2329));
    CascadeMux I__272 (
            .O(N__2354),
            .I(N__2326));
    CascadeMux I__271 (
            .O(N__2353),
            .I(N__2323));
    CascadeMux I__270 (
            .O(N__2352),
            .I(N__2320));
    CascadeMux I__269 (
            .O(N__2351),
            .I(N__2317));
    CascadeMux I__268 (
            .O(N__2350),
            .I(N__2314));
    CascadeMux I__267 (
            .O(N__2349),
            .I(N__2311));
    CascadeMux I__266 (
            .O(N__2348),
            .I(N__2308));
    CascadeMux I__265 (
            .O(N__2347),
            .I(N__2305));
    CascadeMux I__264 (
            .O(N__2346),
            .I(N__2302));
    CascadeMux I__263 (
            .O(N__2345),
            .I(N__2299));
    CascadeMux I__262 (
            .O(N__2344),
            .I(N__2296));
    InMux I__261 (
            .O(N__2341),
            .I(N__2280));
    InMux I__260 (
            .O(N__2338),
            .I(N__2280));
    InMux I__259 (
            .O(N__2335),
            .I(N__2280));
    InMux I__258 (
            .O(N__2332),
            .I(N__2280));
    InMux I__257 (
            .O(N__2329),
            .I(N__2271));
    InMux I__256 (
            .O(N__2326),
            .I(N__2271));
    InMux I__255 (
            .O(N__2323),
            .I(N__2271));
    InMux I__254 (
            .O(N__2320),
            .I(N__2271));
    InMux I__253 (
            .O(N__2317),
            .I(N__2262));
    InMux I__252 (
            .O(N__2314),
            .I(N__2262));
    InMux I__251 (
            .O(N__2311),
            .I(N__2262));
    InMux I__250 (
            .O(N__2308),
            .I(N__2262));
    InMux I__249 (
            .O(N__2305),
            .I(N__2253));
    InMux I__248 (
            .O(N__2302),
            .I(N__2253));
    InMux I__247 (
            .O(N__2299),
            .I(N__2253));
    InMux I__246 (
            .O(N__2296),
            .I(N__2253));
    CascadeMux I__245 (
            .O(N__2295),
            .I(N__2250));
    CascadeMux I__244 (
            .O(N__2294),
            .I(N__2247));
    CascadeMux I__243 (
            .O(N__2293),
            .I(N__2244));
    CascadeMux I__242 (
            .O(N__2292),
            .I(N__2241));
    CascadeMux I__241 (
            .O(N__2291),
            .I(N__2238));
    CascadeMux I__240 (
            .O(N__2290),
            .I(N__2235));
    CascadeMux I__239 (
            .O(N__2289),
            .I(N__2232));
    LocalMux I__238 (
            .O(N__2280),
            .I(N__2227));
    LocalMux I__237 (
            .O(N__2271),
            .I(N__2227));
    LocalMux I__236 (
            .O(N__2262),
            .I(N__2222));
    LocalMux I__235 (
            .O(N__2253),
            .I(N__2222));
    InMux I__234 (
            .O(N__2250),
            .I(N__2215));
    InMux I__233 (
            .O(N__2247),
            .I(N__2215));
    InMux I__232 (
            .O(N__2244),
            .I(N__2215));
    InMux I__231 (
            .O(N__2241),
            .I(N__2206));
    InMux I__230 (
            .O(N__2238),
            .I(N__2206));
    InMux I__229 (
            .O(N__2235),
            .I(N__2206));
    InMux I__228 (
            .O(N__2232),
            .I(N__2206));
    Odrv12 I__227 (
            .O(N__2227),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__226 (
            .O(N__2222),
            .I(CONSTANT_ONE_NET));
    LocalMux I__225 (
            .O(N__2215),
            .I(CONSTANT_ONE_NET));
    LocalMux I__224 (
            .O(N__2206),
            .I(CONSTANT_ONE_NET));
    InMux I__223 (
            .O(N__2197),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1 ));
    InMux I__222 (
            .O(N__2194),
            .I(bfn_26_21_0_));
    CascadeMux I__221 (
            .O(N__2191),
            .I(un1_M_count_q_axbxc7_m4_0_a2_2_cascade_));
    InMux I__220 (
            .O(N__2188),
            .I(N__2185));
    LocalMux I__219 (
            .O(N__2185),
            .I(N__2182));
    Odrv4 I__218 (
            .O(N__2182),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_CO ));
    InMux I__217 (
            .O(N__2179),
            .I(N__2175));
    InMux I__216 (
            .O(N__2178),
            .I(N__2172));
    LocalMux I__215 (
            .O(N__2175),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_0 ));
    LocalMux I__214 (
            .O(N__2172),
            .I(\sr_chain.M_sr_rest_cycles_qZ0Z_0 ));
    InMux I__213 (
            .O(N__2167),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1 ));
    InMux I__212 (
            .O(N__2164),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1 ));
    InMux I__211 (
            .O(N__2161),
            .I(bfn_26_20_0_));
    InMux I__210 (
            .O(N__2158),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1 ));
    InMux I__209 (
            .O(N__2155),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1 ));
    InMux I__208 (
            .O(N__2152),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1 ));
    InMux I__207 (
            .O(N__2149),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1 ));
    InMux I__206 (
            .O(N__2146),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1 ));
    InMux I__205 (
            .O(N__2143),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1 ));
    InMux I__204 (
            .O(N__2140),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1 ));
    InMux I__203 (
            .O(N__2137),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1 ));
    InMux I__202 (
            .O(N__2134),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1 ));
    InMux I__201 (
            .O(N__2131),
            .I(bfn_26_19_0_));
    InMux I__200 (
            .O(N__2128),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1 ));
    InMux I__199 (
            .O(N__2125),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1 ));
    InMux I__198 (
            .O(N__2122),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1 ));
    InMux I__197 (
            .O(N__2119),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1 ));
    InMux I__196 (
            .O(N__2116),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1 ));
    InMux I__195 (
            .O(N__2113),
            .I(N__2110));
    LocalMux I__194 (
            .O(N__2110),
            .I(\reset_cond.M_stage_qZ0Z_1 ));
    InMux I__193 (
            .O(N__2107),
            .I(N__2104));
    LocalMux I__192 (
            .O(N__2104),
            .I(\reset_cond.M_stage_qZ0Z_0 ));
    InMux I__191 (
            .O(N__2101),
            .I(N__2089));
    InMux I__190 (
            .O(N__2100),
            .I(N__2089));
    InMux I__189 (
            .O(N__2099),
            .I(N__2089));
    InMux I__188 (
            .O(N__2098),
            .I(N__2089));
    LocalMux I__187 (
            .O(N__2089),
            .I(N__2086));
    Span12Mux_v I__186 (
            .O(N__2086),
            .I(N__2083));
    Odrv12 I__185 (
            .O(N__2083),
            .I(rst_n_c));
    InMux I__184 (
            .O(N__2080),
            .I(N__2077));
    LocalMux I__183 (
            .O(N__2077),
            .I(\reset_cond.M_stage_qZ0Z_2 ));
    InMux I__182 (
            .O(N__2074),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1 ));
    InMux I__181 (
            .O(N__2071),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1 ));
    InMux I__180 (
            .O(N__2068),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1 ));
    InMux I__179 (
            .O(N__2065),
            .I(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1 ));
    defparam IN_MUX_bfv_28_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_28_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_28_17_0_));
    defparam IN_MUX_bfv_29_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_29_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_29_18_0_));
    defparam IN_MUX_bfv_26_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_18_0_));
    defparam IN_MUX_bfv_26_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_19_0_ (
            .carryinitin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1 ),
            .carryinitout(bfn_26_19_0_));
    defparam IN_MUX_bfv_26_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_20_0_ (
            .carryinitin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1 ),
            .carryinitout(bfn_26_20_0_));
    defparam IN_MUX_bfv_26_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_21_0_ (
            .carryinitin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1 ),
            .carryinitout(bfn_26_21_0_));
    defparam IN_MUX_bfv_30_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_30_15_0_));
    defparam IN_MUX_bfv_30_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_16_0_ (
            .carryinitin(\sr_chain.un1_M_main_clock_count_q_1_cry_7 ),
            .carryinitout(bfn_30_16_0_));
    defparam IN_MUX_bfv_30_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_17_0_ (
            .carryinitin(\sr_chain.un1_M_main_clock_count_q_1_cry_15 ),
            .carryinitout(bfn_30_17_0_));
    defparam IN_MUX_bfv_30_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_18_0_ (
            .carryinitin(\sr_chain.un1_M_main_clock_count_q_1_cry_23 ),
            .carryinitout(bfn_30_18_0_));
    ICE_GB \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_0  (
            .USERSIGNALTOGLOBALBUFFER(N__3700),
            .GLOBALBUFFEROUTPUT(\sr_chain.N_44_g ));
    ICE_GB \reset_cond.M_stage_q_RNIFG9D_3  (
            .USERSIGNALTOGLOBALBUFFER(N__4696),
            .GLOBALBUFFEROUTPUT(N_108_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \reset_cond.M_stage_q_1_LC_17_13_1 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_1_LC_17_13_1 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_1_LC_17_13_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \reset_cond.M_stage_q_1_LC_17_13_1  (
            .in0(N__2099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2107),
            .lcout(\reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4745),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_2_LC_17_13_2 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_2_LC_17_13_2 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_2_LC_17_13_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \reset_cond.M_stage_q_2_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__2100),
            .in2(_gnd_net_),
            .in3(N__2113),
            .lcout(\reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4745),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_0_LC_17_13_5 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_0_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_0_LC_17_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \reset_cond.M_stage_q_0_LC_17_13_5  (
            .in0(N__2098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4745),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_3_LC_17_13_6 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_3_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_3_LC_17_13_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \reset_cond.M_stage_q_3_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__2101),
            .in2(_gnd_net_),
            .in3(N__2080),
            .lcout(M_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4745),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_26_17_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_26_17_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_26_17_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_26_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_rest_cycles_q_0_LC_26_18_0 .C_ON=1'b1;
    defparam \sr_chain.M_sr_rest_cycles_q_0_LC_26_18_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_0_LC_26_18_0 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_0_LC_26_18_0  (
            .in0(N__4949),
            .in1(N__2179),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_26_18_0_),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1 ),
            .clk(N__4750),
            .ce(),
            .sr(N__3454));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_LUT4_0_LC_26_18_1 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_LUT4_0_LC_26_18_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_LUT4_0_LC_26_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_LUT4_0_LC_26_18_1  (
            .in0(_gnd_net_),
            .in1(N__2529),
            .in2(N__2289),
            .in3(N__2074),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_LUT4_0_LC_26_18_2 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_LUT4_0_LC_26_18_2 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_LUT4_0_LC_26_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_LUT4_0_LC_26_18_2  (
            .in0(_gnd_net_),
            .in1(N__2504),
            .in2(N__2293),
            .in3(N__2071),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_LUT4_0_LC_26_18_3 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_LUT4_0_LC_26_18_3 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_LUT4_0_LC_26_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_LUT4_0_LC_26_18_3  (
            .in0(_gnd_net_),
            .in1(N__2479),
            .in2(N__2290),
            .in3(N__2068),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_LUT4_0_LC_26_18_4 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_LUT4_0_LC_26_18_4 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_LUT4_0_LC_26_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_LUT4_0_LC_26_18_4  (
            .in0(_gnd_net_),
            .in1(N__2374),
            .in2(N__2294),
            .in3(N__2065),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_LUT4_0_LC_26_18_5 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_LUT4_0_LC_26_18_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_LUT4_0_LC_26_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_LUT4_0_LC_26_18_5  (
            .in0(_gnd_net_),
            .in1(N__2657),
            .in2(N__2291),
            .in3(N__2140),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_LUT4_0_LC_26_18_6 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_LUT4_0_LC_26_18_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_LUT4_0_LC_26_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_LUT4_0_LC_26_18_6  (
            .in0(_gnd_net_),
            .in1(N__2562),
            .in2(N__2295),
            .in3(N__2137),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_LUT4_0_LC_26_18_7 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_LUT4_0_LC_26_18_7 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_LUT4_0_LC_26_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_LUT4_0_LC_26_18_7  (
            .in0(_gnd_net_),
            .in1(N__2730),
            .in2(N__2292),
            .in3(N__2134),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_LUT4_0_LC_26_19_0 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_LUT4_0_LC_26_19_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_LUT4_0_LC_26_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_LUT4_0_LC_26_19_0  (
            .in0(_gnd_net_),
            .in1(N__2401),
            .in2(N__2350),
            .in3(N__2131),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_CO ),
            .ltout(),
            .carryin(bfn_26_19_0_),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_LUT4_0_LC_26_19_1 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_LUT4_0_LC_26_19_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_LUT4_0_LC_26_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_LUT4_0_LC_26_19_1  (
            .in0(_gnd_net_),
            .in1(N__2434),
            .in2(N__2347),
            .in3(N__2128),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_LUT4_0_LC_26_19_2 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_LUT4_0_LC_26_19_2 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_LUT4_0_LC_26_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_LUT4_0_LC_26_19_2  (
            .in0(_gnd_net_),
            .in1(N__2455),
            .in2(N__2351),
            .in3(N__2125),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_LUT4_0_LC_26_19_3 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_LUT4_0_LC_26_19_3 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_LUT4_0_LC_26_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_LUT4_0_LC_26_19_3  (
            .in0(_gnd_net_),
            .in1(N__2616),
            .in2(N__2344),
            .in3(N__2122),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_LUT4_0_LC_26_19_4 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_LUT4_0_LC_26_19_4 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_LUT4_0_LC_26_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_LUT4_0_LC_26_19_4  (
            .in0(_gnd_net_),
            .in1(N__3222),
            .in2(N__2348),
            .in3(N__2119),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_LUT4_0_LC_26_19_5 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_LUT4_0_LC_26_19_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_LUT4_0_LC_26_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_LUT4_0_LC_26_19_5  (
            .in0(_gnd_net_),
            .in1(N__3198),
            .in2(N__2345),
            .in3(N__2116),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_LUT4_0_LC_26_19_6 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_LUT4_0_LC_26_19_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_LUT4_0_LC_26_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_LUT4_0_LC_26_19_6  (
            .in0(_gnd_net_),
            .in1(N__3176),
            .in2(N__2349),
            .in3(N__2167),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_LUT4_0_LC_26_19_7 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_LUT4_0_LC_26_19_7 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_LUT4_0_LC_26_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_LUT4_0_LC_26_19_7  (
            .in0(_gnd_net_),
            .in1(N__3136),
            .in2(N__2346),
            .in3(N__2164),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_LUT4_0_LC_26_20_0 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_LUT4_0_LC_26_20_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_LUT4_0_LC_26_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_LUT4_0_LC_26_20_0  (
            .in0(_gnd_net_),
            .in1(N__3082),
            .in2(N__2352),
            .in3(N__2161),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_CO ),
            .ltout(),
            .carryin(bfn_26_20_0_),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_LUT4_0_LC_26_20_1 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_LUT4_0_LC_26_20_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_LUT4_0_LC_26_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_LUT4_0_LC_26_20_1  (
            .in0(_gnd_net_),
            .in1(N__3099),
            .in2(N__2356),
            .in3(N__2158),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_LUT4_0_LC_26_20_2 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_LUT4_0_LC_26_20_2 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_LUT4_0_LC_26_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_LUT4_0_LC_26_20_2  (
            .in0(_gnd_net_),
            .in1(N__3059),
            .in2(N__2353),
            .in3(N__2155),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_LUT4_0_LC_26_20_3 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_LUT4_0_LC_26_20_3 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_LUT4_0_LC_26_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_LUT4_0_LC_26_20_3  (
            .in0(_gnd_net_),
            .in1(N__3039),
            .in2(N__2357),
            .in3(N__2152),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_LUT4_0_LC_26_20_4 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_LUT4_0_LC_26_20_4 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_LUT4_0_LC_26_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_LUT4_0_LC_26_20_4  (
            .in0(_gnd_net_),
            .in1(N__3517),
            .in2(N__2354),
            .in3(N__2149),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_LUT4_0_LC_26_20_5 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_LUT4_0_LC_26_20_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_LUT4_0_LC_26_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_LUT4_0_LC_26_20_5  (
            .in0(_gnd_net_),
            .in1(N__3481),
            .in2(N__2358),
            .in3(N__2146),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_LUT4_0_LC_26_20_6 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_LUT4_0_LC_26_20_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_LUT4_0_LC_26_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_LUT4_0_LC_26_20_6  (
            .in0(_gnd_net_),
            .in1(N__3550),
            .in2(N__2355),
            .in3(N__2143),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_LUT4_0_LC_26_20_7 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_LUT4_0_LC_26_20_7 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_LUT4_0_LC_26_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_LUT4_0_LC_26_20_7  (
            .in0(_gnd_net_),
            .in1(N__3012),
            .in2(N__2359),
            .in3(N__2197),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_CO ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_LUT4_0_LC_26_21_0 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_LUT4_0_LC_26_21_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_LUT4_0_LC_26_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_LUT4_0_LC_26_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2194),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNO_1_7_LC_27_14_4.C_ON=1'b0;
    defparam M_count_q_RNO_1_7_LC_27_14_4.SEQ_MODE=4'b0000;
    defparam M_count_q_RNO_1_7_LC_27_14_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_count_q_RNO_1_7_LC_27_14_4 (
            .in0(N__3368),
            .in1(N__3421),
            .in2(N__3324),
            .in3(N__2770),
            .lcout(),
            .ltout(un1_M_count_q_axbxc7_m4_0_a2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNO_0_7_LC_27_14_5.C_ON=1'b0;
    defparam M_count_q_RNO_0_7_LC_27_14_5.SEQ_MODE=4'b0000;
    defparam M_count_q_RNO_0_7_LC_27_14_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_count_q_RNO_0_7_LC_27_14_5 (
            .in0(N__2977),
            .in1(N__2911),
            .in2(N__2191),
            .in3(N__2941),
            .lcout(un1_M_count_q_axbxc7_m4_0_a2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_1_LC_27_15_0.C_ON=1'b0;
    defparam M_count_q_1_LC_27_15_0.SEQ_MODE=4'b1000;
    defparam M_count_q_1_LC_27_15_0.LUT_INIT=16'b1100011011001100;
    LogicCell40 M_count_q_1_LC_27_15_0 (
            .in0(N__4951),
            .in1(N__3425),
            .in2(N__4531),
            .in3(N__2773),
            .lcout(M_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4746),
            .ce(),
            .sr(N__4694));
    defparam M_count_q_3_LC_27_15_4.C_ON=1'b0;
    defparam M_count_q_3_LC_27_15_4.SEQ_MODE=4'b1000;
    defparam M_count_q_3_LC_27_15_4.LUT_INIT=16'b0101111110100000;
    LogicCell40 M_count_q_3_LC_27_15_4 (
            .in0(N__2955),
            .in1(_gnd_net_),
            .in2(N__3380),
            .in3(N__3320),
            .lcout(M_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4746),
            .ce(),
            .sr(N__4694));
    defparam M_count_q_2_LC_27_15_5.C_ON=1'b0;
    defparam M_count_q_2_LC_27_15_5.SEQ_MODE=4'b1000;
    defparam M_count_q_2_LC_27_15_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_count_q_2_LC_27_15_5 (
            .in0(_gnd_net_),
            .in1(N__3370),
            .in2(_gnd_net_),
            .in3(N__2954),
            .lcout(M_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4746),
            .ce(),
            .sr(N__4694));
    defparam M_count_q_0_LC_27_15_7.C_ON=1'b0;
    defparam M_count_q_0_LC_27_15_7.SEQ_MODE=4'b1000;
    defparam M_count_q_0_LC_27_15_7.LUT_INIT=16'b1001100110101010;
    LogicCell40 M_count_q_0_LC_27_15_7 (
            .in0(N__2772),
            .in1(N__4524),
            .in2(_gnd_net_),
            .in3(N__4952),
            .lcout(M_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4746),
            .ce(),
            .sr(N__4694));
    defparam \sr_chain.M_sr_rest_cycles_q_9_LC_27_16_2 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_9_LC_27_16_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_9_LC_27_16_2 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_9_LC_27_16_2  (
            .in0(N__2188),
            .in1(N__3628),
            .in2(_gnd_net_),
            .in3(N__2433),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4748),
            .ce(),
            .sr(N__3460));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_RNO_LC_27_17_0 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_RNO_LC_27_17_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_RNO_LC_27_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_RNO_LC_27_17_0  (
            .in0(N__2528),
            .in1(N__2178),
            .in2(N__2505),
            .in3(N__2477),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_1_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_rest_cycles_q_1_LC_27_17_1 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_1_LC_27_17_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_1_LC_27_17_1 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_1_LC_27_17_1  (
            .in0(N__2530),
            .in1(N__2536),
            .in2(_gnd_net_),
            .in3(N__3617),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4751),
            .ce(),
            .sr(N__3458));
    defparam \sr_chain.M_sr_rest_cycles_q_2_LC_27_17_2 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_2_LC_27_17_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_2_LC_27_17_2 .LUT_INIT=16'b1101001011010010;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_2_LC_27_17_2  (
            .in0(N__3618),
            .in1(N__2512),
            .in2(N__2506),
            .in3(_gnd_net_),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4751),
            .ce(),
            .sr(N__3458));
    defparam \sr_chain.M_sr_rest_cycles_q_3_LC_27_17_3 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_3_LC_27_17_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_3_LC_27_17_3 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_3_LC_27_17_3  (
            .in0(N__2478),
            .in1(N__2485),
            .in2(_gnd_net_),
            .in3(N__3619),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4751),
            .ce(),
            .sr(N__3458));
    defparam \sr_chain.M_sr_rest_cycles_q_10_LC_27_17_4 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_10_LC_27_17_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_10_LC_27_17_4 .LUT_INIT=16'b1100110000111100;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_10_LC_27_17_4  (
            .in0(_gnd_net_),
            .in1(N__2450),
            .in2(N__3626),
            .in3(N__2464),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4751),
            .ce(),
            .sr(N__3458));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_RNO_LC_27_17_5 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_RNO_LC_27_17_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_RNO_LC_27_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_RNO_LC_27_17_5  (
            .in0(N__2396),
            .in1(N__2615),
            .in2(N__2454),
            .in3(N__2429),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_1_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_rest_cycles_q_8_LC_27_17_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_8_LC_27_17_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_8_LC_27_17_6 .LUT_INIT=16'b1100110000111100;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_8_LC_27_17_6  (
            .in0(_gnd_net_),
            .in1(N__2397),
            .in2(N__3627),
            .in3(N__2413),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4751),
            .ce(),
            .sr(N__3458));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_RNO_LC_27_18_0 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_RNO_LC_27_18_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_RNO_LC_27_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_RNO_LC_27_18_0  (
            .in0(N__2561),
            .in1(N__2729),
            .in2(N__2658),
            .in3(N__2372),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_1_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_rest_cycles_q_4_LC_27_18_1 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_4_LC_27_18_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_4_LC_27_18_1 .LUT_INIT=16'b1010010110101010;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_4_LC_27_18_1  (
            .in0(N__2373),
            .in1(_gnd_net_),
            .in2(N__2383),
            .in3(N__3598),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4755),
            .ce(),
            .sr(N__3457));
    defparam \sr_chain.M_sr_rest_cycles_q_5_LC_27_18_2 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_5_LC_27_18_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_5_LC_27_18_2 .LUT_INIT=16'b1101001011010010;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_5_LC_27_18_2  (
            .in0(N__3599),
            .in1(N__2665),
            .in2(N__2659),
            .in3(_gnd_net_),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4755),
            .ce(),
            .sr(N__3457));
    defparam \sr_chain.M_sr_rest_cycles_q_24_LC_27_18_5 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_24_LC_27_18_5 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_24_LC_27_18_5 .LUT_INIT=16'b1111101010001101;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_24_LC_27_18_5  (
            .in0(N__4940),
            .in1(N__4122),
            .in2(N__2638),
            .in3(N__3250),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4755),
            .ce(),
            .sr(N__3457));
    defparam \sr_chain.M_sr_rest_cycles_q_11_LC_27_18_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_11_LC_27_18_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_11_LC_27_18_6 .LUT_INIT=16'b1110111011000011;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_11_LC_27_18_6  (
            .in0(N__4120),
            .in1(N__2617),
            .in2(N__2626),
            .in3(N__4941),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4755),
            .ce(),
            .sr(N__3457));
    defparam \sr_chain.M_sr_rest_cycles_q_12_LC_27_18_7 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_12_LC_27_18_7 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_12_LC_27_18_7 .LUT_INIT=16'b1111100010101101;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_12_LC_27_18_7  (
            .in0(N__4939),
            .in1(N__4121),
            .in2(N__3226),
            .in3(N__2599),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4755),
            .ce(),
            .sr(N__3457));
    defparam \sr_chain.M_sr_rest_cycles_q_13_LC_27_19_0 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_13_LC_27_19_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_13_LC_27_19_0 .LUT_INIT=16'b1111101011000011;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_13_LC_27_19_0  (
            .in0(N__4105),
            .in1(N__2593),
            .in2(N__3205),
            .in3(N__4936),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4758),
            .ce(),
            .sr(N__3455));
    defparam \sr_chain.M_sr_rest_cycles_q_14_LC_27_19_1 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_14_LC_27_19_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_14_LC_27_19_1 .LUT_INIT=16'b1111100010101101;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_14_LC_27_19_1  (
            .in0(N__4934),
            .in1(N__4106),
            .in2(N__3181),
            .in3(N__2587),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4758),
            .ce(),
            .sr(N__3455));
    defparam \sr_chain.M_sr_rest_cycles_q_17_LC_27_19_3 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_17_LC_27_19_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_17_LC_27_19_3 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_17_LC_27_19_3  (
            .in0(N__2581),
            .in1(N__3595),
            .in2(_gnd_net_),
            .in3(N__3100),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4758),
            .ce(),
            .sr(N__3455));
    defparam \sr_chain.M_sr_rest_cycles_q_6_LC_27_19_4 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_6_LC_27_19_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_6_LC_27_19_4 .LUT_INIT=16'b1110111011000011;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_6_LC_27_19_4  (
            .in0(N__4109),
            .in1(N__2563),
            .in2(N__2575),
            .in3(N__4938),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4758),
            .ce(),
            .sr(N__3455));
    defparam \sr_chain.M_sr_rest_cycles_q_19_LC_27_19_5 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_19_LC_27_19_5 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_19_LC_27_19_5 .LUT_INIT=16'b1111101010001101;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_19_LC_27_19_5  (
            .in0(N__4935),
            .in1(N__4108),
            .in2(N__2545),
            .in3(N__3040),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4758),
            .ce(),
            .sr(N__3455));
    defparam \sr_chain.M_sr_rest_cycles_q_18_LC_27_19_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_18_LC_27_19_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_18_LC_27_19_6 .LUT_INIT=16'b1110111011000011;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_18_LC_27_19_6  (
            .in0(N__4107),
            .in1(N__3060),
            .in2(N__2746),
            .in3(N__4937),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4758),
            .ce(),
            .sr(N__3455));
    defparam \sr_chain.M_sr_rest_cycles_q_7_LC_27_19_7 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_7_LC_27_19_7 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_7_LC_27_19_7 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_7_LC_27_19_7  (
            .in0(N__2737),
            .in1(N__3596),
            .in2(_gnd_net_),
            .in3(N__2731),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4758),
            .ce(),
            .sr(N__3455));
    defparam \sr_chain.M_sr_rest_cycles_q_23_LC_27_20_7 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_23_LC_27_20_7 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_23_LC_27_20_7 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_23_LC_27_20_7  (
            .in0(N__2713),
            .in1(N__3597),
            .in2(_gnd_net_),
            .in3(N__3013),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4761),
            .ce(),
            .sr(N__3453));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIH9O82_LC_27_21_5 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIH9O82_LC_27_21_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIH9O82_LC_27_21_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIH9O82_LC_27_21_5  (
            .in0(_gnd_net_),
            .in1(N__4950),
            .in2(_gnd_net_),
            .in3(N__4123),
            .lcout(sr_chain_latch_e1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_7_LC_28_14_1.C_ON=1'b0;
    defparam M_count_q_7_LC_28_14_1.SEQ_MODE=4'b1000;
    defparam M_count_q_7_LC_28_14_1.LUT_INIT=16'b1100011011001100;
    LogicCell40 M_count_q_7_LC_28_14_1 (
            .in0(N__4932),
            .in1(N__2677),
            .in2(N__4510),
            .in3(N__2683),
            .lcout(M_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4747),
            .ce(),
            .sr(N__4695));
    defparam M_count_q_RNIR63U_7_LC_28_14_2.C_ON=1'b0;
    defparam M_count_q_RNIR63U_7_LC_28_14_2.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIR63U_7_LC_28_14_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 M_count_q_RNIR63U_7_LC_28_14_2 (
            .in0(N__2785),
            .in1(N__2676),
            .in2(_gnd_net_),
            .in3(N__3286),
            .lcout(sr_data_to_send_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIQ53U_6_LC_28_14_3.C_ON=1'b0;
    defparam M_count_q_RNIQ53U_6_LC_28_14_3.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIQ53U_6_LC_28_14_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 M_count_q_RNIQ53U_6_LC_28_14_3 (
            .in0(N__3285),
            .in1(N__2976),
            .in2(_gnd_net_),
            .in3(N__2797),
            .lcout(sr_data_to_send_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIO33U_4_LC_28_14_4.C_ON=1'b0;
    defparam M_count_q_RNIO33U_4_LC_28_14_4.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIO33U_4_LC_28_14_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 M_count_q_RNIO33U_4_LC_28_14_4 (
            .in0(N__2940),
            .in1(N__3283),
            .in2(_gnd_net_),
            .in3(N__2842),
            .lcout(sr_data_to_send_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIP43U_5_LC_28_14_5.C_ON=1'b0;
    defparam M_count_q_RNIP43U_5_LC_28_14_5.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIP43U_5_LC_28_14_5.LUT_INIT=16'b1101100011011000;
    LogicCell40 M_count_q_RNIP43U_5_LC_28_14_5 (
            .in0(N__3284),
            .in1(N__2910),
            .in2(N__2821),
            .in3(_gnd_net_),
            .lcout(sr_data_to_send_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_is_sending_q_RNI73BG_0_LC_28_14_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_is_sending_q_RNI73BG_0_LC_28_14_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_is_sending_q_RNI73BG_0_LC_28_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \sr_chain.M_sr_is_sending_q_RNI73BG_0_LC_28_14_6  (
            .in0(_gnd_net_),
            .in1(N__4493),
            .in2(_gnd_net_),
            .in3(N__4931),
            .lcout(sr_chain_is_sending_0_clk),
            .ltout(sr_chain_is_sending_0_clk_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIKV2U_0_LC_28_14_7.C_ON=1'b0;
    defparam M_count_q_RNIKV2U_0_LC_28_14_7.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIKV2U_0_LC_28_14_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 M_count_q_RNIKV2U_0_LC_28_14_7 (
            .in0(_gnd_net_),
            .in1(N__2771),
            .in2(N__2863),
            .in3(N__3657),
            .lcout(sr_data_to_send_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_data_buffer_q_esr_1_LC_28_15_0 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_esr_1_LC_28_15_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_esr_1_LC_28_15_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_esr_1_LC_28_15_0  (
            .in0(N__3639),
            .in1(N__3396),
            .in2(_gnd_net_),
            .in3(N__4484),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4749),
            .ce(N__3670),
            .sr(N__4693));
    defparam \sr_chain.M_sr_data_buffer_q_esr_2_LC_28_15_1 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_esr_2_LC_28_15_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_esr_2_LC_28_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_esr_2_LC_28_15_1  (
            .in0(N__3336),
            .in1(N__2860),
            .in2(_gnd_net_),
            .in3(N__4530),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4749),
            .ce(N__3670),
            .sr(N__4693));
    defparam \sr_chain.M_sr_data_buffer_q_esr_3_LC_28_15_2 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_esr_3_LC_28_15_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_esr_3_LC_28_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_esr_3_LC_28_15_2  (
            .in0(N__3261),
            .in1(N__2854),
            .in2(_gnd_net_),
            .in3(N__4485),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4749),
            .ce(N__3670),
            .sr(N__4693));
    defparam \sr_chain.M_sr_data_buffer_q_esr_4_LC_28_15_3 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_esr_4_LC_28_15_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_esr_4_LC_28_15_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_esr_4_LC_28_15_3  (
            .in0(N__2848),
            .in1(N__4528),
            .in2(_gnd_net_),
            .in3(N__2841),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4749),
            .ce(N__3670),
            .sr(N__4693));
    defparam \sr_chain.M_sr_data_buffer_q_esr_5_LC_28_15_4 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_esr_5_LC_28_15_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_esr_5_LC_28_15_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_esr_5_LC_28_15_4  (
            .in0(N__2830),
            .in1(N__4482),
            .in2(_gnd_net_),
            .in3(N__2817),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4749),
            .ce(N__3670),
            .sr(N__4693));
    defparam \sr_chain.M_sr_data_buffer_q_esr_6_LC_28_15_5 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_esr_6_LC_28_15_5 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_esr_6_LC_28_15_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_esr_6_LC_28_15_5  (
            .in0(N__2806),
            .in1(N__4529),
            .in2(_gnd_net_),
            .in3(N__2796),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4749),
            .ce(N__3670),
            .sr(N__4693));
    defparam \sr_chain.M_sr_data_buffer_q_esr_7_LC_28_15_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_esr_7_LC_28_15_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_esr_7_LC_28_15_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_esr_7_LC_28_15_6  (
            .in0(N__4587),
            .in1(N__4483),
            .in2(_gnd_net_),
            .in3(N__2784),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4749),
            .ce(N__3670),
            .sr(N__4693));
    defparam M_count_q_RNI2TQB1_1_LC_28_16_1.C_ON=1'b0;
    defparam M_count_q_RNI2TQB1_1_LC_28_16_1.SEQ_MODE=4'b0000;
    defparam M_count_q_RNI2TQB1_1_LC_28_16_1.LUT_INIT=16'b0010000000000000;
    LogicCell40 M_count_q_RNI2TQB1_1_LC_28_16_1 (
            .in0(N__2769),
            .in1(N__4479),
            .in2(N__3426),
            .in3(N__4881),
            .lcout(un1_M_count_q_c2),
            .ltout(un1_M_count_q_c2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIIR2L2_4_LC_28_16_2.C_ON=1'b0;
    defparam M_count_q_RNIIR2L2_4_LC_28_16_2.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIIR2L2_4_LC_28_16_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_count_q_RNIIR2L2_4_LC_28_16_2 (
            .in0(N__2932),
            .in1(N__3318),
            .in2(N__2983),
            .in3(N__3369),
            .lcout(un1_M_count_q_c5),
            .ltout(un1_M_count_q_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_6_LC_28_16_3.C_ON=1'b0;
    defparam M_count_q_6_LC_28_16_3.SEQ_MODE=4'b1000;
    defparam M_count_q_6_LC_28_16_3.LUT_INIT=16'b0011111111000000;
    LogicCell40 M_count_q_6_LC_28_16_3 (
            .in0(_gnd_net_),
            .in1(N__2909),
            .in2(N__2980),
            .in3(N__2975),
            .lcout(M_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4752),
            .ce(),
            .sr(N__4692));
    defparam M_count_q_4_LC_28_16_4.C_ON=1'b0;
    defparam M_count_q_4_LC_28_16_4.SEQ_MODE=4'b1000;
    defparam M_count_q_4_LC_28_16_4.LUT_INIT=16'b0110101010101010;
    LogicCell40 M_count_q_4_LC_28_16_4 (
            .in0(N__2933),
            .in1(N__3319),
            .in2(N__3385),
            .in3(N__2956),
            .lcout(M_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4752),
            .ce(),
            .sr(N__4692));
    defparam M_count_q_5_LC_28_16_5.C_ON=1'b0;
    defparam M_count_q_5_LC_28_16_5.SEQ_MODE=4'b1000;
    defparam M_count_q_5_LC_28_16_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_count_q_5_LC_28_16_5 (
            .in0(_gnd_net_),
            .in1(N__2908),
            .in2(_gnd_net_),
            .in3(N__2917),
            .lcout(M_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4752),
            .ce(),
            .sr(N__4692));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_LC_28_17_0 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_LC_28_17_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_LC_28_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_LC_28_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2884),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_28_17_0_),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_LC_28_17_1 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_LC_28_17_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_LC_28_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_LC_28_17_1  (
            .in0(_gnd_net_),
            .in1(N__2875),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_1_0 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_1_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_LC_28_17_2 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_LC_28_17_2 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_LC_28_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_LC_28_17_2  (
            .in0(_gnd_net_),
            .in1(N__2869),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_1_1 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_1_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_LC_28_17_3 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_LC_28_17_3 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_LC_28_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_LC_28_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3157),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_1_2 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_1_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_LC_28_17_4 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_LC_28_17_4 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_LC_28_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_LC_28_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3022),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_1_3 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_1_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_LC_28_17_5 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_LC_28_17_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_LC_28_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_LC_28_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2995),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_1_4 ),
            .carryout(\sr_chain.un1_M_sr_rest_cycles_q_1_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_inv_LC_28_17_6 .C_ON=1'b1;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_inv_LC_28_17_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_inv_LC_28_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_inv_LC_28_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3238),
            .in3(N__3249),
            .lcout(\sr_chain.M_sr_rest_cycles_q_i_24 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_sr_rest_cycles_q_1_5 ),
            .carryout(sr_chain_un1_M_sr_rest_cycles_q_1_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_LUT4_0_LC_28_17_7.C_ON=1'b0;
    defparam sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_LUT4_0_LC_28_17_7.SEQ_MODE=4'b0000;
    defparam sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_LUT4_0_LC_28_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_LUT4_0_LC_28_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3229),
            .lcout(sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_RNO_LC_28_18_0 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_RNO_LC_28_18_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_RNO_LC_28_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_RNO_LC_28_18_0  (
            .in0(N__3221),
            .in1(N__3197),
            .in2(N__3180),
            .in3(N__3128),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_1_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_rest_cycles_q_15_LC_28_18_1 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_15_LC_28_18_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_15_LC_28_18_1 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_15_LC_28_18_1  (
            .in0(N__3129),
            .in1(N__3148),
            .in2(_gnd_net_),
            .in3(N__3594),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4759),
            .ce(),
            .sr(N__3459));
    defparam \sr_chain.M_sr_rest_cycles_q_16_LC_28_18_4 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_16_LC_28_18_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_16_LC_28_18_4 .LUT_INIT=16'b1110111010100101;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_16_LC_28_18_4  (
            .in0(N__3075),
            .in1(N__4101),
            .in2(N__3115),
            .in3(N__4907),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4759),
            .ce(),
            .sr(N__3459));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_RNO_LC_28_18_5 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_RNO_LC_28_18_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_RNO_LC_28_18_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_RNO_LC_28_18_5  (
            .in0(N__3098),
            .in1(N__3074),
            .in2(N__3061),
            .in3(N__3038),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_1_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_RNO_LC_28_19_0 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_RNO_LC_28_19_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_RNO_LC_28_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_RNO_LC_28_19_0  (
            .in0(N__3545),
            .in1(N__3476),
            .in2(N__3516),
            .in3(N__3011),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_1_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIFAS5_LC_28_19_6 .C_ON=1'b0;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIFAS5_LC_28_19_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIFAS5_LC_28_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIFAS5_LC_28_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4933),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_1_6_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_rest_cycles_q_22_LC_28_20_2 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_22_LC_28_20_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_22_LC_28_20_2 .LUT_INIT=16'b1110111011000011;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_22_LC_28_20_2  (
            .in0(N__4104),
            .in1(N__3549),
            .in2(N__3562),
            .in3(N__4944),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4763),
            .ce(),
            .sr(N__3456));
    defparam \sr_chain.M_sr_rest_cycles_q_20_LC_28_20_4 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_20_LC_28_20_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_20_LC_28_20_4 .LUT_INIT=16'b1110111011000011;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_20_LC_28_20_4  (
            .in0(N__4102),
            .in1(N__3515),
            .in2(N__3529),
            .in3(N__4942),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4763),
            .ce(),
            .sr(N__3456));
    defparam \sr_chain.M_sr_rest_cycles_q_21_LC_28_20_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_rest_cycles_q_21_LC_28_20_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_rest_cycles_q_21_LC_28_20_6 .LUT_INIT=16'b1110111011000011;
    LogicCell40 \sr_chain.M_sr_rest_cycles_q_21_LC_28_20_6  (
            .in0(N__4103),
            .in1(N__3480),
            .in2(N__3493),
            .in3(N__4943),
            .lcout(\sr_chain.M_sr_rest_cycles_qZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4763),
            .ce(),
            .sr(N__3456));
    defparam M_count_q_RNIL03U_1_LC_29_14_1.C_ON=1'b0;
    defparam M_count_q_RNIL03U_1_LC_29_14_1.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIL03U_1_LC_29_14_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 M_count_q_RNIL03U_1_LC_29_14_1 (
            .in0(N__3397),
            .in1(N__3430),
            .in2(_gnd_net_),
            .in3(N__3287),
            .lcout(sr_data_to_send_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIM13U_2_LC_29_14_4.C_ON=1'b0;
    defparam M_count_q_RNIM13U_2_LC_29_14_4.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIM13U_2_LC_29_14_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 M_count_q_RNIM13U_2_LC_29_14_4 (
            .in0(N__3288),
            .in1(N__3384),
            .in2(_gnd_net_),
            .in3(N__3337),
            .lcout(sr_data_to_send_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_count_q_RNIN23U_3_LC_29_14_5.C_ON=1'b0;
    defparam M_count_q_RNIN23U_3_LC_29_14_5.SEQ_MODE=4'b0000;
    defparam M_count_q_RNIN23U_3_LC_29_14_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 M_count_q_RNIN23U_3_LC_29_14_5 (
            .in0(N__3325),
            .in1(N__3289),
            .in2(_gnd_net_),
            .in3(N__3262),
            .lcout(sr_data_to_send_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_4_c_RNO_LC_29_15_0 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_4_c_RNO_LC_29_15_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_4_c_RNO_LC_29_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.M_main_clock_count_d8_4_c_RNO_LC_29_15_0  (
            .in0(N__4236),
            .in1(N__4200),
            .in2(N__4258),
            .in3(N__4185),
            .lcout(\sr_chain.M_main_clock_count_d8_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_RNIL1D81_1_LC_29_15_1 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_RNIL1D81_1_LC_29_15_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_clock_count_q_RNIL1D81_1_LC_29_15_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \sr_chain.M_sr_clock_count_q_RNIL1D81_1_LC_29_15_1  (
            .in0(N__4008),
            .in1(_gnd_net_),
            .in2(N__3688),
            .in3(N__3716),
            .lcout(\sr_chain.un1_M_sr_clock_count_q_1_c2 ),
            .ltout(\sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_2_LC_29_15_2 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_2_LC_29_15_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_clock_count_q_2_LC_29_15_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \sr_chain.M_sr_clock_count_q_2_LC_29_15_2  (
            .in0(N__3884),
            .in1(_gnd_net_),
            .in2(N__3691),
            .in3(N__3932),
            .lcout(\sr_chain.M_sr_clock_count_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4753),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_3_c_RNO_LC_29_15_3 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_3_c_RNO_LC_29_15_3 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_3_c_RNO_LC_29_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.M_main_clock_count_d8_3_c_RNO_LC_29_15_3  (
            .in0(N__3847),
            .in1(N__4272),
            .in2(N__3832),
            .in3(N__3813),
            .lcout(\sr_chain.M_main_clock_count_d8_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_1_LC_29_15_4 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_1_LC_29_15_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_clock_count_q_1_LC_29_15_4 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \sr_chain.M_sr_clock_count_q_1_LC_29_15_4  (
            .in0(N__3718),
            .in1(N__3687),
            .in2(N__3888),
            .in3(N__4010),
            .lcout(\sr_chain.M_sr_clock_count_qZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4753),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_RNI74IL_3_LC_29_15_5 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_RNI74IL_3_LC_29_15_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_clock_count_q_RNI74IL_3_LC_29_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \sr_chain.M_sr_clock_count_q_RNI74IL_3_LC_29_15_5  (
            .in0(N__3931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3902),
            .lcout(),
            .ltout(\sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_RNIV7TL1_1_LC_29_15_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_RNIV7TL1_1_LC_29_15_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_clock_count_q_RNIV7TL1_1_LC_29_15_6 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \sr_chain.M_sr_clock_count_q_RNIV7TL1_1_LC_29_15_6  (
            .in0(N__3950),
            .in1(N__3683),
            .in2(N__3673),
            .in3(N__4007),
            .lcout(\sr_chain.un1_M_sr_clock_count_q ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_0_LC_29_15_7 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_0_LC_29_15_7 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_clock_count_q_0_LC_29_15_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \sr_chain.M_sr_clock_count_q_0_LC_29_15_7  (
            .in0(N__4009),
            .in1(N__3880),
            .in2(_gnd_net_),
            .in3(N__3717),
            .lcout(\sr_chain.M_sr_clock_count_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4753),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNIIHTA1_LC_29_16_1 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNIIHTA1_LC_29_16_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNIIHTA1_LC_29_16_1 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \sr_chain.M_main_clock_count_d8_6_c_RNIIHTA1_LC_29_16_1  (
            .in0(N__4662),
            .in1(N__3726),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_data_buffer_q_0_LC_29_16_3 .C_ON=1'b0;
    defparam \sr_chain.M_sr_data_buffer_q_0_LC_29_16_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_data_buffer_q_0_LC_29_16_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \sr_chain.M_sr_data_buffer_q_0_LC_29_16_3  (
            .in0(N__4480),
            .in1(N__3727),
            .in2(N__3643),
            .in3(N__3658),
            .lcout(\sr_chain.M_sr_data_buffer_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4756),
            .ce(),
            .sr(N__4684));
    defparam \sr_chain.M_sr_is_sending_q_LC_29_16_4 .C_ON=1'b0;
    defparam \sr_chain.M_sr_is_sending_q_LC_29_16_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_is_sending_q_LC_29_16_4 .LUT_INIT=16'b1110011011101110;
    LogicCell40 \sr_chain.M_sr_is_sending_q_LC_29_16_4  (
            .in0(N__4854),
            .in1(N__4481),
            .in2(N__4573),
            .in3(N__4060),
            .lcout(sr_chain_latch13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4756),
            .ce(),
            .sr(N__4684));
    defparam \sr_chain.M_sr_is_sending_q_RNI73BG_LC_29_16_5 .C_ON=1'b0;
    defparam \sr_chain.M_sr_is_sending_q_RNI73BG_LC_29_16_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_is_sending_q_RNI73BG_LC_29_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \sr_chain.M_sr_is_sending_q_RNI73BG_LC_29_16_5  (
            .in0(_gnd_net_),
            .in1(N__4454),
            .in2(_gnd_net_),
            .in3(N__4853),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI31KT_LC_29_17_0 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI31KT_LC_29_17_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI31KT_LC_29_17_0 .LUT_INIT=16'b1101010100000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_6_c_RNI31KT_LC_29_17_0  (
            .in0(N__4486),
            .in1(N__4059),
            .in2(N__4027),
            .in3(N__4914),
            .lcout(\sr_chain.un1_M_sr_rest_cycles_q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_1_c_RNO_LC_29_17_1 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_1_c_RNO_LC_29_17_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_1_c_RNO_LC_29_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_1_c_RNO_LC_29_17_1  (
            .in0(N__4332),
            .in1(N__4302),
            .in2(N__4366),
            .in3(N__4287),
            .lcout(\sr_chain.M_main_clock_count_d8_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_is_sending_q_RNIMJKT_LC_29_17_2 .C_ON=1'b0;
    defparam \sr_chain.M_sr_is_sending_q_RNIMJKT_LC_29_17_2 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_is_sending_q_RNIMJKT_LC_29_17_2 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \sr_chain.M_sr_is_sending_q_RNIMJKT_LC_29_17_2  (
            .in0(N__4661),
            .in1(_gnd_net_),
            .in2(N__4509),
            .in3(N__4916),
            .lcout(\sr_chain.M_sr_is_sending_q_RNIMJKTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_0_c_RNO_LC_29_17_3 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_0_c_RNO_LC_29_17_3 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_0_c_RNO_LC_29_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_0_c_RNO_LC_29_17_3  (
            .in0(N__4380),
            .in1(N__4137),
            .in2(N__4222),
            .in3(N__4395),
            .lcout(\sr_chain.M_main_clock_count_d8_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNII1RI_LC_29_17_4 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNII1RI_LC_29_17_4 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNII1RI_LC_29_17_4 .LUT_INIT=16'b1100110000001100;
    LogicCell40 \sr_chain.M_main_clock_count_d8_6_c_RNII1RI_LC_29_17_4  (
            .in0(_gnd_net_),
            .in1(N__4915),
            .in2(N__4508),
            .in3(N__4058),
            .lcout(\sr_chain.M_main_clock_count_d_0_sqmuxa ),
            .ltout(\sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_LC_29_17_5 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_LC_29_17_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_LC_29_17_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_LC_29_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3703),
            .in3(N__4660),
            .lcout(\sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_5_c_RNO_LC_29_17_6 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_5_c_RNO_LC_29_17_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_5_c_RNO_LC_29_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sr_chain.M_main_clock_count_d8_5_c_RNO_LC_29_17_6  (
            .in0(N__4317),
            .in1(N__4347),
            .in2(N__4171),
            .in3(N__4152),
            .lcout(\sr_chain.M_main_clock_count_d8_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_2_c_RNO_LC_29_17_7 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_2_c_RNO_LC_29_17_7 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_2_c_RNO_LC_29_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_2_c_RNO_LC_29_17_7  (
            .in0(N__5059),
            .in1(N__4989),
            .in2(N__5026),
            .in3(N__5040),
            .lcout(\sr_chain.M_main_clock_count_d8_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_0_c_LC_29_18_0 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_d8_0_c_LC_29_18_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_0_c_LC_29_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_0_c_LC_29_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3799),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_29_18_0_),
            .carryout(\sr_chain.M_main_clock_count_d8_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_1_c_LC_29_18_1 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_d8_1_c_LC_29_18_1 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_1_c_LC_29_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_1_c_LC_29_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3790),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.M_main_clock_count_d8_0 ),
            .carryout(\sr_chain.M_main_clock_count_d8_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_2_c_LC_29_18_2 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_d8_2_c_LC_29_18_2 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_2_c_LC_29_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_2_c_LC_29_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3781),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.M_main_clock_count_d8_1 ),
            .carryout(\sr_chain.M_main_clock_count_d8_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_3_c_LC_29_18_3 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_d8_3_c_LC_29_18_3 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_3_c_LC_29_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_3_c_LC_29_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.M_main_clock_count_d8_2 ),
            .carryout(\sr_chain.M_main_clock_count_d8_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_4_c_LC_29_18_4 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_d8_4_c_LC_29_18_4 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_4_c_LC_29_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_4_c_LC_29_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3760),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.M_main_clock_count_d8_3 ),
            .carryout(\sr_chain.M_main_clock_count_d8_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_5_c_LC_29_18_5 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_d8_5_c_LC_29_18_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_5_c_LC_29_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_5_c_LC_29_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\sr_chain.M_main_clock_count_d8_4 ),
            .carryout(\sr_chain.M_main_clock_count_d8_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_6_c_inv_LC_29_18_6 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_d8_6_c_inv_LC_29_18_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_6_c_inv_LC_29_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sr_chain.M_main_clock_count_d8_6_c_inv_LC_29_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3739),
            .in3(N__5007),
            .lcout(\sr_chain.M_main_clock_count_q_i_23 ),
            .ltout(),
            .carryin(\sr_chain.M_main_clock_count_d8_5 ),
            .carryout(\sr_chain.M_main_clock_count_d8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_THRU_LUT4_0_LC_29_18_7 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_THRU_LUT4_0_LC_29_18_7 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_THRU_LUT4_0_LC_29_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_THRU_LUT4_0_LC_29_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3730),
            .lcout(\sr_chain.M_main_clock_count_d8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_bit_q_RNO_0_LC_29_19_0 .C_ON=1'b0;
    defparam \sr_chain.M_sr_bit_q_RNO_0_LC_29_19_0 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_bit_q_RNO_0_LC_29_19_0 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \sr_chain.M_sr_bit_q_RNO_0_LC_29_19_0  (
            .in0(N__4022),
            .in1(N__4498),
            .in2(N__3964),
            .in3(N__4053),
            .lcout(\sr_chain.M_sr_bit_d_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI2VR22_LC_29_19_4 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI2VR22_LC_29_19_4 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNI2VR22_LC_29_19_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_6_c_RNI2VR22_LC_29_19_4  (
            .in0(N__4570),
            .in1(N__4497),
            .in2(_gnd_net_),
            .in3(N__4052),
            .lcout(\sr_chain.latch_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNIPG9U1_LC_29_19_5 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNIPG9U1_LC_29_19_5 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_main_clock_count_d8_6_c_RNIPG9U1_LC_29_19_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \sr_chain.M_main_clock_count_d8_6_c_RNIPG9U1_LC_29_19_5  (
            .in0(N__4054),
            .in1(N__4571),
            .in2(_gnd_net_),
            .in3(N__4945),
            .lcout(),
            .ltout(\sr_chain.M_sr_bit_d12_m_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_RNIHJDP2_0_LC_29_19_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_RNIHJDP2_0_LC_29_19_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_clock_count_q_RNIHJDP2_0_LC_29_19_6 .LUT_INIT=16'b1010111100110011;
    LogicCell40 \sr_chain.M_sr_clock_count_q_RNIHJDP2_0_LC_29_19_6  (
            .in0(N__4023),
            .in1(N__4954),
            .in2(N__3985),
            .in3(N__4499),
            .lcout(sr_clk_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sr_chain.M_sr_clock_count_q_4_LC_30_14_0 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_4_LC_30_14_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_clock_count_q_4_LC_30_14_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \sr_chain.M_sr_clock_count_q_4_LC_30_14_0  (
            .in0(N__3913),
            .in1(N__3904),
            .in2(N__3960),
            .in3(N__3934),
            .lcout(\sr_chain.M_sr_clock_count_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4754),
            .ce(),
            .sr(N__3889));
    defparam \sr_chain.M_sr_clock_count_q_3_LC_30_14_1 .C_ON=1'b0;
    defparam \sr_chain.M_sr_clock_count_q_3_LC_30_14_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_clock_count_q_3_LC_30_14_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \sr_chain.M_sr_clock_count_q_3_LC_30_14_1  (
            .in0(N__3903),
            .in1(N__3933),
            .in2(_gnd_net_),
            .in3(N__3912),
            .lcout(\sr_chain.M_sr_clock_count_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4754),
            .ce(),
            .sr(N__3889));
    defparam \sr_chain.M_main_clock_count_q_0_LC_30_15_0 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_0_LC_30_15_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_0_LC_30_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_0_LC_30_15_0  (
            .in0(_gnd_net_),
            .in1(N__3846),
            .in2(N__3862),
            .in3(N__3861),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_30_15_0_),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_0 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_1_LC_30_15_1 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_1_LC_30_15_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_1_LC_30_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_1_LC_30_15_1  (
            .in0(_gnd_net_),
            .in1(N__3831),
            .in2(_gnd_net_),
            .in3(N__3817),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_1 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_0 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_1 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_2_LC_30_15_2 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_2_LC_30_15_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_2_LC_30_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_2_LC_30_15_2  (
            .in0(_gnd_net_),
            .in1(N__3814),
            .in2(_gnd_net_),
            .in3(N__3802),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_2 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_1 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_2 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_3_LC_30_15_3 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_3_LC_30_15_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_3_LC_30_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_3_LC_30_15_3  (
            .in0(_gnd_net_),
            .in1(N__4273),
            .in2(_gnd_net_),
            .in3(N__4261),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_3 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_2 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_3 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_4_LC_30_15_4 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_4_LC_30_15_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_4_LC_30_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_4_LC_30_15_4  (
            .in0(_gnd_net_),
            .in1(N__4254),
            .in2(_gnd_net_),
            .in3(N__4240),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_4 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_3 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_4 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_5_LC_30_15_5 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_5_LC_30_15_5 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_5_LC_30_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_5_LC_30_15_5  (
            .in0(_gnd_net_),
            .in1(N__4237),
            .in2(_gnd_net_),
            .in3(N__4225),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_5 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_4 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_5 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_6_LC_30_15_6 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_6_LC_30_15_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_6_LC_30_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_6_LC_30_15_6  (
            .in0(_gnd_net_),
            .in1(N__4218),
            .in2(_gnd_net_),
            .in3(N__4204),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_6 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_5 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_6 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_7_LC_30_15_7 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_7_LC_30_15_7 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_7_LC_30_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_7_LC_30_15_7  (
            .in0(_gnd_net_),
            .in1(N__4201),
            .in2(_gnd_net_),
            .in3(N__4189),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_7 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_6 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_7 ),
            .clk(N__4757),
            .ce(),
            .sr(N__4978));
    defparam \sr_chain.M_main_clock_count_q_8_LC_30_16_0 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_8_LC_30_16_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_8_LC_30_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_8_LC_30_16_0  (
            .in0(_gnd_net_),
            .in1(N__4186),
            .in2(_gnd_net_),
            .in3(N__4174),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_8 ),
            .ltout(),
            .carryin(bfn_30_16_0_),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_8 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_9_LC_30_16_1 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_9_LC_30_16_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_9_LC_30_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_9_LC_30_16_1  (
            .in0(_gnd_net_),
            .in1(N__4170),
            .in2(_gnd_net_),
            .in3(N__4156),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_9 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_8 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_9 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_10_LC_30_16_2 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_10_LC_30_16_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_10_LC_30_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_10_LC_30_16_2  (
            .in0(_gnd_net_),
            .in1(N__4153),
            .in2(_gnd_net_),
            .in3(N__4141),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_10 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_9 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_10 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_11_LC_30_16_3 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_11_LC_30_16_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_11_LC_30_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_11_LC_30_16_3  (
            .in0(_gnd_net_),
            .in1(N__4138),
            .in2(_gnd_net_),
            .in3(N__4126),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_11 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_10 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_11 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_12_LC_30_16_4 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_12_LC_30_16_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_12_LC_30_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_12_LC_30_16_4  (
            .in0(_gnd_net_),
            .in1(N__4396),
            .in2(_gnd_net_),
            .in3(N__4384),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_12 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_11 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_12 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_13_LC_30_16_5 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_13_LC_30_16_5 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_13_LC_30_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_13_LC_30_16_5  (
            .in0(_gnd_net_),
            .in1(N__4381),
            .in2(_gnd_net_),
            .in3(N__4369),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_13 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_12 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_13 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_14_LC_30_16_6 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_14_LC_30_16_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_14_LC_30_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_14_LC_30_16_6  (
            .in0(_gnd_net_),
            .in1(N__4365),
            .in2(_gnd_net_),
            .in3(N__4351),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_14 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_13 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_14 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_15_LC_30_16_7 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_15_LC_30_16_7 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_15_LC_30_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_15_LC_30_16_7  (
            .in0(_gnd_net_),
            .in1(N__4348),
            .in2(_gnd_net_),
            .in3(N__4336),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_15 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_14 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_15 ),
            .clk(N__4760),
            .ce(),
            .sr(N__4976));
    defparam \sr_chain.M_main_clock_count_q_16_LC_30_17_0 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_16_LC_30_17_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_16_LC_30_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_16_LC_30_17_0  (
            .in0(_gnd_net_),
            .in1(N__4333),
            .in2(_gnd_net_),
            .in3(N__4321),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_16 ),
            .ltout(),
            .carryin(bfn_30_17_0_),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_16 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_17_LC_30_17_1 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_17_LC_30_17_1 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_17_LC_30_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_17_LC_30_17_1  (
            .in0(_gnd_net_),
            .in1(N__4318),
            .in2(_gnd_net_),
            .in3(N__4306),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_17 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_16 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_17 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_18_LC_30_17_2 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_18_LC_30_17_2 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_18_LC_30_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_18_LC_30_17_2  (
            .in0(_gnd_net_),
            .in1(N__4303),
            .in2(_gnd_net_),
            .in3(N__4291),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_18 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_17 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_18 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_19_LC_30_17_3 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_19_LC_30_17_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_19_LC_30_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_19_LC_30_17_3  (
            .in0(_gnd_net_),
            .in1(N__4288),
            .in2(_gnd_net_),
            .in3(N__4276),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_19 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_18 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_19 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_20_LC_30_17_4 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_20_LC_30_17_4 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_20_LC_30_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_20_LC_30_17_4  (
            .in0(_gnd_net_),
            .in1(N__5058),
            .in2(_gnd_net_),
            .in3(N__5044),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_20 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_19 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_20 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_21_LC_30_17_5 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_21_LC_30_17_5 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_21_LC_30_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_21_LC_30_17_5  (
            .in0(_gnd_net_),
            .in1(N__5041),
            .in2(_gnd_net_),
            .in3(N__5029),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_21 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_20 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_21 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_22_LC_30_17_6 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_22_LC_30_17_6 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_22_LC_30_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_22_LC_30_17_6  (
            .in0(_gnd_net_),
            .in1(N__5025),
            .in2(_gnd_net_),
            .in3(N__5011),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_22 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_21 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_22 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_23_LC_30_17_7 .C_ON=1'b1;
    defparam \sr_chain.M_main_clock_count_q_23_LC_30_17_7 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_23_LC_30_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sr_chain.M_main_clock_count_q_23_LC_30_17_7  (
            .in0(_gnd_net_),
            .in1(N__5008),
            .in2(_gnd_net_),
            .in3(N__4996),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_23 ),
            .ltout(),
            .carryin(\sr_chain.un1_M_main_clock_count_q_1_cry_22 ),
            .carryout(\sr_chain.un1_M_main_clock_count_q_1_cry_23 ),
            .clk(N__4762),
            .ce(),
            .sr(N__4975));
    defparam \sr_chain.M_main_clock_count_q_24_LC_30_18_0 .C_ON=1'b0;
    defparam \sr_chain.M_main_clock_count_q_24_LC_30_18_0 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_main_clock_count_q_24_LC_30_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \sr_chain.M_main_clock_count_q_24_LC_30_18_0  (
            .in0(_gnd_net_),
            .in1(N__4990),
            .in2(_gnd_net_),
            .in3(N__4993),
            .lcout(\sr_chain.M_main_clock_count_qZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4764),
            .ce(),
            .sr(N__4977));
    defparam \sr_chain.M_sr_bit_q_LC_30_19_3 .C_ON=1'b0;
    defparam \sr_chain.M_sr_bit_q_LC_30_19_3 .SEQ_MODE=4'b1000;
    defparam \sr_chain.M_sr_bit_q_LC_30_19_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \sr_chain.M_sr_bit_q_LC_30_19_3  (
            .in0(N__4408),
            .in1(N__4960),
            .in2(N__4782),
            .in3(N__4953),
            .lcout(sr_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4765),
            .ce(),
            .sr(N__4688));
    defparam \sr_chain.M_sr_bit_q_RNO_1_LC_31_15_6 .C_ON=1'b0;
    defparam \sr_chain.M_sr_bit_q_RNO_1_LC_31_15_6 .SEQ_MODE=4'b0000;
    defparam \sr_chain.M_sr_bit_q_RNO_1_LC_31_15_6 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \sr_chain.M_sr_bit_q_RNO_1_LC_31_15_6  (
            .in0(N__4588),
            .in1(N__4572),
            .in2(N__4543),
            .in3(N__4511),
            .lcout(\sr_chain.M_sr_bit_q_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
