-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Oct 30 2022 12:29:41

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    sr_latch : out std_logic;
    sr_data : out std_logic;
    sr_clk : out std_logic;
    rst_n : in std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2182\ : std_logic;
signal \N__2179\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2172\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2125\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2065\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal rst_n_c : std_logic;
signal \reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \bfn_26_18_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1\ : std_logic;
signal \bfn_26_19_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1\ : std_logic;
signal \bfn_26_20_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1\ : std_logic;
signal \bfn_26_21_0_\ : std_logic;
signal \un1_M_count_q_axbxc7_m4_0_a2_2_cascade_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_0\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_2\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_3\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_10\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_9\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_8\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_4\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_5\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_11\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_6\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_7\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_CO\ : std_logic;
signal sr_chain_latch_e1_i : std_logic;
signal \un1_M_count_q_axbxc7_m4_0_a2_3\ : std_logic;
signal \M_count_qZ0Z_7\ : std_logic;
signal \sr_chain_is_sending_0_clk_cascade_\ : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_1\ : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_2\ : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_3\ : std_logic;
signal sr_data_to_send_4 : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_4\ : std_logic;
signal sr_data_to_send_5 : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_5\ : std_logic;
signal sr_data_to_send_6 : std_logic;
signal sr_data_to_send_7 : std_logic;
signal \M_count_qZ0Z_0\ : std_logic;
signal \un1_M_count_q_c2_cascade_\ : std_logic;
signal \un1_M_count_q_c5_cascade_\ : std_logic;
signal \M_count_qZ0Z_6\ : std_logic;
signal \un1_M_count_q_c2\ : std_logic;
signal \M_count_qZ0Z_4\ : std_logic;
signal \un1_M_count_q_c5\ : std_logic;
signal \M_count_qZ0Z_5\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_0_and\ : std_logic;
signal \bfn_28_17_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_1_and\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_0\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_2_and\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_2\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_3\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_4\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_24\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_q_i_24\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_5\ : std_logic;
signal \sr_chain_un1_M_sr_rest_cycles_q_1_6\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_12\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_13\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_14\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_3_and\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_15\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_17\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_16\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_18\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_19\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_4_and\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_23\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_5_and\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_22\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_20\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_21\ : std_logic;
signal \N_108_g\ : std_logic;
signal \M_count_qZ0Z_1\ : std_logic;
signal sr_data_to_send_1 : std_logic;
signal \M_count_qZ0Z_2\ : std_logic;
signal sr_data_to_send_2 : std_logic;
signal \M_count_qZ0Z_3\ : std_logic;
signal sr_chain_is_sending_0_clk : std_logic;
signal sr_data_to_send_3 : std_logic;
signal \sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ1Z_1\ : std_logic;
signal \sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_5_0_0\ : std_logic;
signal sr_data_to_send_0 : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_0\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_5_0\ : std_logic;
signal \sr_chain.M_main_clock_count_d_0_sqmuxa\ : std_logic;
signal \sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_0_and\ : std_logic;
signal \bfn_29_18_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_1_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_0\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_2_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_1\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_3_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_2\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_4_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_3\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_5_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_4\ : std_logic;
signal \sr_chain.M_main_clock_count_q_i_23\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_5\ : std_logic;
signal \sr_chain.M_main_clock_count_d8\ : std_logic;
signal \sr_chain.latch_0_sqmuxa_1\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_0\ : std_logic;
signal \sr_chain.M_sr_bit_d12_m_0_cascade_\ : std_logic;
signal sr_clk_c : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_4\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_2\ : std_logic;
signal \sr_chain.un1_M_sr_clock_count_q_1_c2\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_3\ : std_logic;
signal \sr_chain.M_sr_is_sending_q_RNIMJKTZ0\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_3_0\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_0\ : std_logic;
signal \bfn_30_15_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_1\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_0\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_2\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_1\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_3\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_2\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_4\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_3\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_5\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_4\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_6\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_5\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_7\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_6\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_7\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_8\ : std_logic;
signal \bfn_30_16_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_9\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_8\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_10\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_9\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_11\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_10\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_12\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_11\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_13\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_12\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_14\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_13\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_15\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_14\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_15\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_16\ : std_logic;
signal \bfn_30_17_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_17\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_16\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_18\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_17\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_19\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_18\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_20\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_19\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_21\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_20\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_22\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_21\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_23\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_22\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_23\ : std_logic;
signal \bfn_30_18_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_24\ : std_logic;
signal \sr_chain.N_44_g\ : std_logic;
signal \sr_chain.M_sr_bit_d_2_sqmuxa\ : std_logic;
signal \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\ : std_logic;
signal sr_data_c : std_logic;
signal clk_c_g : std_logic;
signal \M_reset_cond_out_0\ : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_6\ : std_logic;
signal \sr_chain.un1_M_sr_clock_count_q\ : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_7\ : std_logic;
signal sr_chain_latch13 : std_logic;
signal \sr_chain.M_sr_bit_q_3\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal rst_n_wire : std_logic;
signal sr_clk_wire : std_logic;
signal sr_data_wire : std_logic;
signal sr_latch_wire : std_logic;

begin
    clk_wire <= clk;
    rst_n_wire <= rst_n;
    sr_clk <= sr_clk_wire;
    sr_data <= sr_data_wire;
    sr_latch <= sr_latch_wire;

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5114\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5116\,
            DIN => \N__5115\,
            DOUT => \N__5114\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5116\,
            PADOUT => \N__5115\,
            PADIN => \N__5114\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5105\,
            DIN => \N__5104\,
            DOUT => \N__5103\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5105\,
            PADOUT => \N__5104\,
            PADIN => \N__5103\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \sr_clk_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5096\,
            DIN => \N__5095\,
            DOUT => \N__5094\,
            PACKAGEPIN => sr_clk_wire
        );

    \sr_clk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5096\,
            PADOUT => \N__5095\,
            PADIN => \N__5094\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3982\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \sr_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5087\,
            DIN => \N__5086\,
            DOUT => \N__5085\,
            PACKAGEPIN => sr_data_wire
        );

    \sr_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5087\,
            PADOUT => \N__5086\,
            PADIN => \N__5085\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4798\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \sr_latch_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5078\,
            DIN => \N__5077\,
            DOUT => \N__5076\,
            PACKAGEPIN => sr_latch_wire
        );

    \sr_latch_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5078\,
            PADOUT => \N__5077\,
            PADIN => \N__5076\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2707\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1177\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5055\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5052\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5052\,
            I => \sr_chain.M_main_clock_count_qZ0Z_20\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__5049\,
            I => \sr_chain.M_main_clock_count_qZ0Z_20\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5044\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_19\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5037\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5034\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5037\,
            I => \sr_chain.M_main_clock_count_qZ0Z_21\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5034\,
            I => \sr_chain.M_main_clock_count_qZ0Z_21\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5029\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_20\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__5026\,
            I => \N__5022\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5019\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5016\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5019\,
            I => \sr_chain.M_main_clock_count_qZ0Z_22\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5016\,
            I => \sr_chain.M_main_clock_count_qZ0Z_22\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5011\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_21\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5004\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5001\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5004\,
            I => \sr_chain.M_main_clock_count_qZ0Z_23\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5001\,
            I => \sr_chain.M_main_clock_count_qZ0Z_23\
        );

    \I__1156\ : InMux
    port map (
            O => \N__4996\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_22\
        );

    \I__1155\ : InMux
    port map (
            O => \N__4993\,
            I => \bfn_30_18_0_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4986\
        );

    \I__1153\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4983\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__4986\,
            I => \sr_chain.M_main_clock_count_qZ0Z_24\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__4983\,
            I => \sr_chain.M_main_clock_count_qZ0Z_24\
        );

    \I__1150\ : SRMux
    port map (
            O => \N__4978\,
            I => \N__4966\
        );

    \I__1149\ : SRMux
    port map (
            O => \N__4977\,
            I => \N__4966\
        );

    \I__1148\ : SRMux
    port map (
            O => \N__4976\,
            I => \N__4966\
        );

    \I__1147\ : SRMux
    port map (
            O => \N__4975\,
            I => \N__4966\
        );

    \I__1146\ : GlobalMux
    port map (
            O => \N__4966\,
            I => \N__4963\
        );

    \I__1145\ : gio2CtrlBuf
    port map (
            O => \N__4963\,
            I => \sr_chain.N_44_g\
        );

    \I__1144\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4957\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__4957\,
            I => \sr_chain.M_sr_bit_d_2_sqmuxa\
        );

    \I__1142\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4946\
        );

    \I__1141\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4928\
        );

    \I__1140\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4923\
        );

    \I__1139\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4923\
        );

    \I__1138\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4920\
        );

    \I__1137\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4917\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__4946\,
            I => \N__4911\
        );

    \I__1135\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4908\
        );

    \I__1134\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4900\
        );

    \I__1133\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4900\
        );

    \I__1132\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4900\
        );

    \I__1131\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4893\
        );

    \I__1130\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4893\
        );

    \I__1129\ : InMux
    port map (
            O => \N__4939\,
            I => \N__4893\
        );

    \I__1128\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4882\
        );

    \I__1127\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4882\
        );

    \I__1126\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4882\
        );

    \I__1125\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4882\
        );

    \I__1124\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4882\
        );

    \I__1123\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4878\
        );

    \I__1122\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4873\
        );

    \I__1121\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4873\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4870\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__4923\,
            I => \N__4867\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4862\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__4917\,
            I => \N__4862\
        );

    \I__1116\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4855\
        );

    \I__1115\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4855\
        );

    \I__1114\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4855\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__4911\,
            I => \N__4850\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4847\
        );

    \I__1111\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4844\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4837\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__4893\,
            I => \N__4837\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__4882\,
            I => \N__4837\
        );

    \I__1107\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4834\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__4878\,
            I => \N__4829\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__4873\,
            I => \N__4829\
        );

    \I__1104\ : Span4Mux_v
    port map (
            O => \N__4870\,
            I => \N__4820\
        );

    \I__1103\ : Span4Mux_v
    port map (
            O => \N__4867\,
            I => \N__4820\
        );

    \I__1102\ : Span4Mux_v
    port map (
            O => \N__4862\,
            I => \N__4820\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__4855\,
            I => \N__4820\
        );

    \I__1100\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4815\
        );

    \I__1099\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4815\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__4850\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1097\ : Odrv4
    port map (
            O => \N__4847\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__4844\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__4837\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__4834\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1093\ : Odrv12
    port map (
            O => \N__4829\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__4820\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4815\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__1090\ : IoInMux
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4795\,
            I => \N__4792\
        );

    \I__1088\ : IoSpan4Mux
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__1087\ : Span4Mux_s2_h
    port map (
            O => \N__4789\,
            I => \N__4786\
        );

    \I__1086\ : Sp12to4
    port map (
            O => \N__4786\,
            I => \N__4783\
        );

    \I__1085\ : Span12Mux_s10_h
    port map (
            O => \N__4783\,
            I => \N__4779\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__4782\,
            I => \N__4776\
        );

    \I__1083\ : Span12Mux_h
    port map (
            O => \N__4779\,
            I => \N__4773\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4770\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__4773\,
            I => sr_data_c
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4770\,
            I => sr_data_c
        );

    \I__1079\ : ClkMux
    port map (
            O => \N__4765\,
            I => \N__4702\
        );

    \I__1078\ : ClkMux
    port map (
            O => \N__4764\,
            I => \N__4702\
        );

    \I__1077\ : ClkMux
    port map (
            O => \N__4763\,
            I => \N__4702\
        );

    \I__1076\ : ClkMux
    port map (
            O => \N__4762\,
            I => \N__4702\
        );

    \I__1075\ : ClkMux
    port map (
            O => \N__4761\,
            I => \N__4702\
        );

    \I__1074\ : ClkMux
    port map (
            O => \N__4760\,
            I => \N__4702\
        );

    \I__1073\ : ClkMux
    port map (
            O => \N__4759\,
            I => \N__4702\
        );

    \I__1072\ : ClkMux
    port map (
            O => \N__4758\,
            I => \N__4702\
        );

    \I__1071\ : ClkMux
    port map (
            O => \N__4757\,
            I => \N__4702\
        );

    \I__1070\ : ClkMux
    port map (
            O => \N__4756\,
            I => \N__4702\
        );

    \I__1069\ : ClkMux
    port map (
            O => \N__4755\,
            I => \N__4702\
        );

    \I__1068\ : ClkMux
    port map (
            O => \N__4754\,
            I => \N__4702\
        );

    \I__1067\ : ClkMux
    port map (
            O => \N__4753\,
            I => \N__4702\
        );

    \I__1066\ : ClkMux
    port map (
            O => \N__4752\,
            I => \N__4702\
        );

    \I__1065\ : ClkMux
    port map (
            O => \N__4751\,
            I => \N__4702\
        );

    \I__1064\ : ClkMux
    port map (
            O => \N__4750\,
            I => \N__4702\
        );

    \I__1063\ : ClkMux
    port map (
            O => \N__4749\,
            I => \N__4702\
        );

    \I__1062\ : ClkMux
    port map (
            O => \N__4748\,
            I => \N__4702\
        );

    \I__1061\ : ClkMux
    port map (
            O => \N__4747\,
            I => \N__4702\
        );

    \I__1060\ : ClkMux
    port map (
            O => \N__4746\,
            I => \N__4702\
        );

    \I__1059\ : ClkMux
    port map (
            O => \N__4745\,
            I => \N__4702\
        );

    \I__1058\ : GlobalMux
    port map (
            O => \N__4702\,
            I => \N__4699\
        );

    \I__1057\ : gio2CtrlBuf
    port map (
            O => \N__4699\,
            I => clk_c_g
        );

    \I__1056\ : IoInMux
    port map (
            O => \N__4696\,
            I => \N__4689\
        );

    \I__1055\ : SRMux
    port map (
            O => \N__4695\,
            I => \N__4685\
        );

    \I__1054\ : SRMux
    port map (
            O => \N__4694\,
            I => \N__4681\
        );

    \I__1053\ : SRMux
    port map (
            O => \N__4693\,
            I => \N__4678\
        );

    \I__1052\ : SRMux
    port map (
            O => \N__4692\,
            I => \N__4675\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4689\,
            I => \N__4672\
        );

    \I__1050\ : SRMux
    port map (
            O => \N__4688\,
            I => \N__4669\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4685\,
            I => \N__4666\
        );

    \I__1048\ : SRMux
    port map (
            O => \N__4684\,
            I => \N__4663\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4655\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__4678\,
            I => \N__4655\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4675\,
            I => \N__4652\
        );

    \I__1044\ : Span4Mux_s1_v
    port map (
            O => \N__4672\,
            I => \N__4649\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__4669\,
            I => \N__4646\
        );

    \I__1042\ : Span4Mux_v
    port map (
            O => \N__4666\,
            I => \N__4641\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4663\,
            I => \N__4641\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4638\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4633\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4633\
        );

    \I__1037\ : Span4Mux_v
    port map (
            O => \N__4655\,
            I => \N__4630\
        );

    \I__1036\ : Span4Mux_v
    port map (
            O => \N__4652\,
            I => \N__4627\
        );

    \I__1035\ : Sp12to4
    port map (
            O => \N__4649\,
            I => \N__4624\
        );

    \I__1034\ : Span4Mux_h
    port map (
            O => \N__4646\,
            I => \N__4621\
        );

    \I__1033\ : Sp12to4
    port map (
            O => \N__4641\,
            I => \N__4614\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4638\,
            I => \N__4614\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4633\,
            I => \N__4614\
        );

    \I__1030\ : Span4Mux_h
    port map (
            O => \N__4630\,
            I => \N__4609\
        );

    \I__1029\ : Span4Mux_h
    port map (
            O => \N__4627\,
            I => \N__4609\
        );

    \I__1028\ : Span12Mux_h
    port map (
            O => \N__4624\,
            I => \N__4606\
        );

    \I__1027\ : Sp12to4
    port map (
            O => \N__4621\,
            I => \N__4601\
        );

    \I__1026\ : Span12Mux_v
    port map (
            O => \N__4614\,
            I => \N__4601\
        );

    \I__1025\ : Span4Mux_h
    port map (
            O => \N__4609\,
            I => \N__4598\
        );

    \I__1024\ : Span12Mux_v
    port map (
            O => \N__4606\,
            I => \N__4593\
        );

    \I__1023\ : Span12Mux_h
    port map (
            O => \N__4601\,
            I => \N__4593\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__4598\,
            I => \M_reset_cond_out_0\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__4593\,
            I => \M_reset_cond_out_0\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4584\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4581\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4584\,
            I => \N__4578\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4581\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_6\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__4578\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_6\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__4573\,
            I => \N__4567\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4564\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4559\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4559\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4567\,
            I => \N__4556\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4564\,
            I => \N__4553\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4559\,
            I => \N__4550\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__4556\,
            I => \sr_chain.un1_M_sr_clock_count_q\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__4553\,
            I => \sr_chain.un1_M_sr_clock_count_q\
        );

    \I__1006\ : Odrv12
    port map (
            O => \N__4550\,
            I => \sr_chain.un1_M_sr_clock_count_q\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__4543\,
            I => \N__4540\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4537\,
            I => \N__4534\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__4534\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_7\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__4531\,
            I => \N__4525\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4517\
        );

    \I__999\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4517\
        );

    \I__998\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4517\
        );

    \I__997\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4512\
        );

    \I__996\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4512\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4503\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4512\,
            I => \N__4503\
        );

    \I__993\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4500\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__4510\,
            I => \N__4494\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__4509\,
            I => \N__4490\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4508\,
            I => \N__4487\
        );

    \I__989\ : Span4Mux_h
    port map (
            O => \N__4503\,
            I => \N__4474\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4500\,
            I => \N__4474\
        );

    \I__987\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4467\
        );

    \I__986\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4467\
        );

    \I__985\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4467\
        );

    \I__984\ : InMux
    port map (
            O => \N__4494\,
            I => \N__4462\
        );

    \I__983\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4462\
        );

    \I__982\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4455\
        );

    \I__981\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4455\
        );

    \I__980\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4455\
        );

    \I__979\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4445\
        );

    \I__978\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4445\
        );

    \I__977\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4445\
        );

    \I__976\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4445\
        );

    \I__975\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4440\
        );

    \I__974\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4440\
        );

    \I__973\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4437\
        );

    \I__972\ : Span4Mux_s3_h
    port map (
            O => \N__4474\,
            I => \N__4432\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4467\,
            I => \N__4432\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4429\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4455\,
            I => \N__4426\
        );

    \I__968\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4423\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4445\,
            I => sr_chain_latch13
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4440\,
            I => sr_chain_latch13
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4437\,
            I => sr_chain_latch13
        );

    \I__964\ : Odrv4
    port map (
            O => \N__4432\,
            I => sr_chain_latch13
        );

    \I__963\ : Odrv4
    port map (
            O => \N__4429\,
            I => sr_chain_latch13
        );

    \I__962\ : Odrv4
    port map (
            O => \N__4426\,
            I => sr_chain_latch13
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4423\,
            I => sr_chain_latch13
        );

    \I__960\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4405\,
            I => \N__4402\
        );

    \I__958\ : Span4Mux_v
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__957\ : Odrv4
    port map (
            O => \N__4399\,
            I => \sr_chain.M_sr_bit_q_3\
        );

    \I__956\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4392\
        );

    \I__955\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4389\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4392\,
            I => \sr_chain.M_main_clock_count_qZ0Z_12\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4389\,
            I => \sr_chain.M_main_clock_count_qZ0Z_12\
        );

    \I__952\ : InMux
    port map (
            O => \N__4384\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_11\
        );

    \I__951\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4377\
        );

    \I__950\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4374\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4377\,
            I => \sr_chain.M_main_clock_count_qZ0Z_13\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4374\,
            I => \sr_chain.M_main_clock_count_qZ0Z_13\
        );

    \I__947\ : InMux
    port map (
            O => \N__4369\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_12\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__4366\,
            I => \N__4362\
        );

    \I__945\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4359\
        );

    \I__944\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4356\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4359\,
            I => \sr_chain.M_main_clock_count_qZ0Z_14\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4356\,
            I => \sr_chain.M_main_clock_count_qZ0Z_14\
        );

    \I__941\ : InMux
    port map (
            O => \N__4351\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_13\
        );

    \I__940\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4344\
        );

    \I__939\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4341\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4344\,
            I => \sr_chain.M_main_clock_count_qZ0Z_15\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4341\,
            I => \sr_chain.M_main_clock_count_qZ0Z_15\
        );

    \I__936\ : InMux
    port map (
            O => \N__4336\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_14\
        );

    \I__935\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4329\
        );

    \I__934\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4326\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4329\,
            I => \sr_chain.M_main_clock_count_qZ0Z_16\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4326\,
            I => \sr_chain.M_main_clock_count_qZ0Z_16\
        );

    \I__931\ : InMux
    port map (
            O => \N__4321\,
            I => \bfn_30_17_0_\
        );

    \I__930\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4314\
        );

    \I__929\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4311\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4314\,
            I => \sr_chain.M_main_clock_count_qZ0Z_17\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4311\,
            I => \sr_chain.M_main_clock_count_qZ0Z_17\
        );

    \I__926\ : InMux
    port map (
            O => \N__4306\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_16\
        );

    \I__925\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4299\
        );

    \I__924\ : InMux
    port map (
            O => \N__4302\,
            I => \N__4296\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4299\,
            I => \sr_chain.M_main_clock_count_qZ0Z_18\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4296\,
            I => \sr_chain.M_main_clock_count_qZ0Z_18\
        );

    \I__921\ : InMux
    port map (
            O => \N__4291\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_17\
        );

    \I__920\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4284\
        );

    \I__919\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4284\,
            I => \sr_chain.M_main_clock_count_qZ0Z_19\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4281\,
            I => \sr_chain.M_main_clock_count_qZ0Z_19\
        );

    \I__916\ : InMux
    port map (
            O => \N__4276\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_18\
        );

    \I__915\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4269\
        );

    \I__914\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4266\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4269\,
            I => \sr_chain.M_main_clock_count_qZ0Z_3\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4266\,
            I => \sr_chain.M_main_clock_count_qZ0Z_3\
        );

    \I__911\ : InMux
    port map (
            O => \N__4261\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_2\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__4258\,
            I => \N__4255\
        );

    \I__909\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4251\
        );

    \I__908\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4248\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4251\,
            I => \N__4245\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4248\,
            I => \sr_chain.M_main_clock_count_qZ0Z_4\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__4245\,
            I => \sr_chain.M_main_clock_count_qZ0Z_4\
        );

    \I__904\ : InMux
    port map (
            O => \N__4240\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_3\
        );

    \I__903\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4233\
        );

    \I__902\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4230\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4233\,
            I => \sr_chain.M_main_clock_count_qZ0Z_5\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4230\,
            I => \sr_chain.M_main_clock_count_qZ0Z_5\
        );

    \I__899\ : InMux
    port map (
            O => \N__4225\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_4\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__897\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4215\
        );

    \I__896\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4212\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4212\,
            I => \sr_chain.M_main_clock_count_qZ0Z_6\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__4209\,
            I => \sr_chain.M_main_clock_count_qZ0Z_6\
        );

    \I__892\ : InMux
    port map (
            O => \N__4204\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_5\
        );

    \I__891\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4197\
        );

    \I__890\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4194\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4197\,
            I => \sr_chain.M_main_clock_count_qZ0Z_7\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4194\,
            I => \sr_chain.M_main_clock_count_qZ0Z_7\
        );

    \I__887\ : InMux
    port map (
            O => \N__4189\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_6\
        );

    \I__886\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4182\
        );

    \I__885\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4179\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4182\,
            I => \sr_chain.M_main_clock_count_qZ0Z_8\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4179\,
            I => \sr_chain.M_main_clock_count_qZ0Z_8\
        );

    \I__882\ : InMux
    port map (
            O => \N__4174\,
            I => \bfn_30_16_0_\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__4171\,
            I => \N__4167\
        );

    \I__880\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4164\
        );

    \I__879\ : InMux
    port map (
            O => \N__4167\,
            I => \N__4161\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4164\,
            I => \sr_chain.M_main_clock_count_qZ0Z_9\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4161\,
            I => \sr_chain.M_main_clock_count_qZ0Z_9\
        );

    \I__876\ : InMux
    port map (
            O => \N__4156\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_8\
        );

    \I__875\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4149\
        );

    \I__874\ : InMux
    port map (
            O => \N__4152\,
            I => \N__4146\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4149\,
            I => \sr_chain.M_main_clock_count_qZ0Z_10\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4146\,
            I => \sr_chain.M_main_clock_count_qZ0Z_10\
        );

    \I__871\ : InMux
    port map (
            O => \N__4141\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_9\
        );

    \I__870\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4134\
        );

    \I__869\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4131\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4134\,
            I => \sr_chain.M_main_clock_count_qZ0Z_11\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4131\,
            I => \sr_chain.M_main_clock_count_qZ0Z_11\
        );

    \I__866\ : InMux
    port map (
            O => \N__4126\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_10\
        );

    \I__865\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4117\
        );

    \I__864\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4110\
        );

    \I__863\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4110\
        );

    \I__862\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4110\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4117\,
            I => \N__4098\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4110\,
            I => \N__4095\
        );

    \I__859\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4084\
        );

    \I__858\ : InMux
    port map (
            O => \N__4108\,
            I => \N__4084\
        );

    \I__857\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4084\
        );

    \I__856\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4084\
        );

    \I__855\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4084\
        );

    \I__854\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4077\
        );

    \I__853\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4077\
        );

    \I__852\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4077\
        );

    \I__851\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4074\
        );

    \I__850\ : Span4Mux_v
    port map (
            O => \N__4098\,
            I => \N__4067\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__4095\,
            I => \N__4067\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4084\,
            I => \N__4067\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4077\,
            I => \sr_chain.latch_0_sqmuxa_1\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4074\,
            I => \sr_chain.latch_0_sqmuxa_1\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__4067\,
            I => \sr_chain.latch_0_sqmuxa_1\
        );

    \I__844\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4055\
        );

    \I__843\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4047\
        );

    \I__842\ : InMux
    port map (
            O => \N__4058\,
            I => \N__4047\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4055\,
            I => \N__4044\
        );

    \I__840\ : InMux
    port map (
            O => \N__4054\,
            I => \N__4037\
        );

    \I__839\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4037\
        );

    \I__838\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4037\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4047\,
            I => \N__4034\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__4044\,
            I => \sr_chain.M_main_clock_count_d8_THRU_CO\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4037\,
            I => \sr_chain.M_main_clock_count_d8_THRU_CO\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__4034\,
            I => \sr_chain.M_main_clock_count_d8_THRU_CO\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__832\ : InMux
    port map (
            O => \N__4024\,
            I => \N__4019\
        );

    \I__831\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4014\
        );

    \I__830\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4014\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4019\,
            I => \N__4011\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4014\,
            I => \N__4004\
        );

    \I__827\ : Span4Mux_s3_h
    port map (
            O => \N__4011\,
            I => \N__4001\
        );

    \I__826\ : InMux
    port map (
            O => \N__4010\,
            I => \N__3992\
        );

    \I__825\ : InMux
    port map (
            O => \N__4009\,
            I => \N__3992\
        );

    \I__824\ : InMux
    port map (
            O => \N__4008\,
            I => \N__3992\
        );

    \I__823\ : InMux
    port map (
            O => \N__4007\,
            I => \N__3992\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__4004\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_0\
        );

    \I__821\ : Odrv4
    port map (
            O => \N__4001\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_0\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__3992\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_0\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__3985\,
            I => \sr_chain.M_sr_bit_d12_m_0_cascade_\
        );

    \I__818\ : IoInMux
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__3979\,
            I => \N__3976\
        );

    \I__816\ : Span12Mux_s4_h
    port map (
            O => \N__3976\,
            I => \N__3973\
        );

    \I__815\ : Span12Mux_h
    port map (
            O => \N__3973\,
            I => \N__3970\
        );

    \I__814\ : Span12Mux_h
    port map (
            O => \N__3970\,
            I => \N__3967\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__3967\,
            I => sr_clk_c
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__3964\,
            I => \N__3961\
        );

    \I__811\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3957\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__3960\,
            I => \N__3954\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__3957\,
            I => \N__3951\
        );

    \I__808\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3947\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__3951\,
            I => \N__3944\
        );

    \I__806\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3941\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3947\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_4\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__3944\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_4\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__3941\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_4\
        );

    \I__802\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3928\
        );

    \I__801\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3925\
        );

    \I__800\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3920\
        );

    \I__799\ : InMux
    port map (
            O => \N__3931\,
            I => \N__3920\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__3928\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_2\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__3925\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_2\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__3920\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_2\
        );

    \I__795\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3907\
        );

    \I__794\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3907\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3907\,
            I => \sr_chain.un1_M_sr_clock_count_q_1_c2\
        );

    \I__792\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3897\
        );

    \I__791\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3897\
        );

    \I__790\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3894\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3897\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_3\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__3894\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_3\
        );

    \I__787\ : SRMux
    port map (
            O => \N__3889\,
            I => \N__3885\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__3888\,
            I => \N__3881\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3885\,
            I => \N__3877\
        );

    \I__784\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3870\
        );

    \I__783\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3870\
        );

    \I__782\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3870\
        );

    \I__781\ : Span4Mux_s3_h
    port map (
            O => \N__3877\,
            I => \N__3865\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__3870\,
            I => \N__3865\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__3865\,
            I => \sr_chain.M_sr_is_sending_q_RNIMJKTZ0\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__3862\,
            I => \N__3858\
        );

    \I__777\ : InMux
    port map (
            O => \N__3861\,
            I => \N__3855\
        );

    \I__776\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3852\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__3855\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_3_0\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3852\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_3_0\
        );

    \I__773\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3843\
        );

    \I__772\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3840\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3843\,
            I => \N__3837\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3840\,
            I => \sr_chain.M_main_clock_count_qZ0Z_0\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__3837\,
            I => \sr_chain.M_main_clock_count_qZ0Z_0\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__3832\,
            I => \N__3828\
        );

    \I__767\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3825\
        );

    \I__766\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3822\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3825\,
            I => \sr_chain.M_main_clock_count_qZ0Z_1\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3822\,
            I => \sr_chain.M_main_clock_count_qZ0Z_1\
        );

    \I__763\ : InMux
    port map (
            O => \N__3817\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_0\
        );

    \I__762\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3810\
        );

    \I__761\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3807\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3810\,
            I => \sr_chain.M_main_clock_count_qZ0Z_2\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3807\,
            I => \sr_chain.M_main_clock_count_qZ0Z_2\
        );

    \I__758\ : InMux
    port map (
            O => \N__3802\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_1\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__3799\,
            I => \N__3796\
        );

    \I__756\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3793\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3793\,
            I => \sr_chain.M_main_clock_count_d8_0_and\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__3790\,
            I => \N__3787\
        );

    \I__753\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3784\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3784\,
            I => \sr_chain.M_main_clock_count_d8_1_and\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__3781\,
            I => \N__3778\
        );

    \I__750\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3775\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3775\,
            I => \sr_chain.M_main_clock_count_d8_2_and\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__3772\,
            I => \N__3769\
        );

    \I__747\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3766\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3766\,
            I => \N__3763\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__3763\,
            I => \sr_chain.M_main_clock_count_d8_3_and\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__3760\,
            I => \N__3757\
        );

    \I__743\ : InMux
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__741\ : Odrv12
    port map (
            O => \N__3751\,
            I => \sr_chain.M_main_clock_count_d8_4_and\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__739\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3742\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3742\,
            I => \sr_chain.M_main_clock_count_d8_5_and\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__3739\,
            I => \N__3736\
        );

    \I__736\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3733\,
            I => \sr_chain.M_main_clock_count_q_i_23\
        );

    \I__734\ : InMux
    port map (
            O => \N__3730\,
            I => \sr_chain.M_main_clock_count_d8\
        );

    \I__733\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3721\
        );

    \I__732\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3721\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3721\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_5_0\
        );

    \I__730\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3709\
        );

    \I__729\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3709\
        );

    \I__728\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3709\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__3706\,
            I => \sr_chain.M_main_clock_count_d_0_sqmuxa\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__3703\,
            I => \sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_\
        );

    \I__724\ : IoInMux
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3697\,
            I => \N__3694\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__3694\,
            I => \sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__3691\,
            I => \sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__3688\,
            I => \N__3684\
        );

    \I__719\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3676\
        );

    \I__718\ : InMux
    port map (
            O => \N__3684\,
            I => \N__3676\
        );

    \I__717\ : InMux
    port map (
            O => \N__3683\,
            I => \N__3676\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3676\,
            I => \sr_chain.M_sr_clock_count_qZ1Z_1\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__3673\,
            I => \sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_\
        );

    \I__714\ : CEMux
    port map (
            O => \N__3670\,
            I => \N__3667\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3667\,
            I => \N__3664\
        );

    \I__712\ : Span4Mux_v
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__3661\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_5_0_0\
        );

    \I__710\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3654\
        );

    \I__709\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3651\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3654\,
            I => \N__3648\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__3651\,
            I => sr_data_to_send_0
        );

    \I__706\ : Odrv4
    port map (
            O => \N__3648\,
            I => sr_data_to_send_0
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__3643\,
            I => \N__3640\
        );

    \I__704\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3636\
        );

    \I__703\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3633\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3636\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_0\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3633\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_0\
        );

    \I__700\ : InMux
    port map (
            O => \N__3628\,
            I => \N__3623\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__3627\,
            I => \N__3620\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__3626\,
            I => \N__3614\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3623\,
            I => \N__3611\
        );

    \I__696\ : InMux
    port map (
            O => \N__3620\,
            I => \N__3600\
        );

    \I__695\ : InMux
    port map (
            O => \N__3619\,
            I => \N__3600\
        );

    \I__694\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3600\
        );

    \I__693\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3600\
        );

    \I__692\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3600\
        );

    \I__691\ : Span4Mux_h
    port map (
            O => \N__3611\,
            I => \N__3589\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3600\,
            I => \N__3589\
        );

    \I__689\ : InMux
    port map (
            O => \N__3599\,
            I => \N__3584\
        );

    \I__688\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3584\
        );

    \I__687\ : InMux
    port map (
            O => \N__3597\,
            I => \N__3581\
        );

    \I__686\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3576\
        );

    \I__685\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3576\
        );

    \I__684\ : InMux
    port map (
            O => \N__3594\,
            I => \N__3573\
        );

    \I__683\ : Odrv4
    port map (
            O => \N__3589\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3584\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3581\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3576\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3573\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__677\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3556\,
            I => \N__3553\
        );

    \I__675\ : Odrv12
    port map (
            O => \N__3553\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_CO\
        );

    \I__674\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3546\
        );

    \I__673\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3542\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3546\,
            I => \N__3539\
        );

    \I__671\ : InMux
    port map (
            O => \N__3545\,
            I => \N__3536\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3542\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_22\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__3539\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_22\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3536\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_22\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__3529\,
            I => \N__3526\
        );

    \I__666\ : InMux
    port map (
            O => \N__3526\,
            I => \N__3523\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3523\,
            I => \N__3520\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__3520\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_CO\
        );

    \I__663\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3512\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__3516\,
            I => \N__3509\
        );

    \I__661\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3506\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3512\,
            I => \N__3503\
        );

    \I__659\ : InMux
    port map (
            O => \N__3509\,
            I => \N__3500\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3506\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_20\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__3503\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_20\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3500\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_20\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__3493\,
            I => \N__3490\
        );

    \I__654\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3487\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__3484\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_CO\
        );

    \I__651\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3477\
        );

    \I__650\ : InMux
    port map (
            O => \N__3480\,
            I => \N__3473\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3477\,
            I => \N__3470\
        );

    \I__648\ : InMux
    port map (
            O => \N__3476\,
            I => \N__3467\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3473\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_21\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__3470\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_21\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3467\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_21\
        );

    \I__644\ : SRMux
    port map (
            O => \N__3460\,
            I => \N__3436\
        );

    \I__643\ : SRMux
    port map (
            O => \N__3459\,
            I => \N__3436\
        );

    \I__642\ : SRMux
    port map (
            O => \N__3458\,
            I => \N__3436\
        );

    \I__641\ : SRMux
    port map (
            O => \N__3457\,
            I => \N__3436\
        );

    \I__640\ : SRMux
    port map (
            O => \N__3456\,
            I => \N__3436\
        );

    \I__639\ : SRMux
    port map (
            O => \N__3455\,
            I => \N__3436\
        );

    \I__638\ : SRMux
    port map (
            O => \N__3454\,
            I => \N__3436\
        );

    \I__637\ : SRMux
    port map (
            O => \N__3453\,
            I => \N__3436\
        );

    \I__636\ : GlobalMux
    port map (
            O => \N__3436\,
            I => \N__3433\
        );

    \I__635\ : gio2CtrlBuf
    port map (
            O => \N__3433\,
            I => \N_108_g\
        );

    \I__634\ : InMux
    port map (
            O => \N__3430\,
            I => \N__3427\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3427\,
            I => \N__3422\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__3426\,
            I => \N__3418\
        );

    \I__631\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3415\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__3422\,
            I => \N__3412\
        );

    \I__629\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3409\
        );

    \I__628\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3406\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3415\,
            I => \M_count_qZ0Z_1\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__3412\,
            I => \M_count_qZ0Z_1\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3409\,
            I => \M_count_qZ0Z_1\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3406\,
            I => \M_count_qZ0Z_1\
        );

    \I__623\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3393\
        );

    \I__622\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3390\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3393\,
            I => sr_data_to_send_1
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3390\,
            I => sr_data_to_send_1
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__3385\,
            I => \N__3381\
        );

    \I__618\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3377\
        );

    \I__617\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3374\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__3380\,
            I => \N__3371\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3377\,
            I => \N__3365\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3374\,
            I => \N__3362\
        );

    \I__613\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3357\
        );

    \I__612\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3357\
        );

    \I__611\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3354\
        );

    \I__610\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3351\
        );

    \I__609\ : Span4Mux_h
    port map (
            O => \N__3365\,
            I => \N__3348\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__3362\,
            I => \M_count_qZ0Z_2\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3357\,
            I => \M_count_qZ0Z_2\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3354\,
            I => \M_count_qZ0Z_2\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3351\,
            I => \M_count_qZ0Z_2\
        );

    \I__604\ : Odrv4
    port map (
            O => \N__3348\,
            I => \M_count_qZ0Z_2\
        );

    \I__603\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3333\
        );

    \I__602\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3330\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3333\,
            I => sr_data_to_send_2
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3330\,
            I => sr_data_to_send_2
        );

    \I__599\ : InMux
    port map (
            O => \N__3325\,
            I => \N__3321\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3324\,
            I => \N__3315\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3321\,
            I => \N__3312\
        );

    \I__596\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3309\
        );

    \I__595\ : InMux
    port map (
            O => \N__3319\,
            I => \N__3304\
        );

    \I__594\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3304\
        );

    \I__593\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3301\
        );

    \I__592\ : Span4Mux_h
    port map (
            O => \N__3312\,
            I => \N__3298\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3309\,
            I => \M_count_qZ0Z_3\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3304\,
            I => \M_count_qZ0Z_3\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3301\,
            I => \M_count_qZ0Z_3\
        );

    \I__588\ : Odrv4
    port map (
            O => \N__3298\,
            I => \M_count_qZ0Z_3\
        );

    \I__587\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3276\
        );

    \I__586\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3276\
        );

    \I__585\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3276\
        );

    \I__584\ : InMux
    port map (
            O => \N__3286\,
            I => \N__3267\
        );

    \I__583\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3267\
        );

    \I__582\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3267\
        );

    \I__581\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3267\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3276\,
            I => sr_chain_is_sending_0_clk
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3267\,
            I => sr_chain_is_sending_0_clk
        );

    \I__578\ : InMux
    port map (
            O => \N__3262\,
            I => \N__3258\
        );

    \I__577\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3255\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3258\,
            I => sr_data_to_send_3
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3255\,
            I => sr_data_to_send_3
        );

    \I__574\ : InMux
    port map (
            O => \N__3250\,
            I => \N__3246\
        );

    \I__573\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3243\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3246\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_24\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3243\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_24\
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__3238\,
            I => \N__3235\
        );

    \I__569\ : InMux
    port map (
            O => \N__3235\,
            I => \N__3232\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3232\,
            I => \sr_chain.M_sr_rest_cycles_q_i_24\
        );

    \I__567\ : InMux
    port map (
            O => \N__3229\,
            I => \sr_chain_un1_M_sr_rest_cycles_q_1_6\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__565\ : InMux
    port map (
            O => \N__3223\,
            I => \N__3218\
        );

    \I__564\ : InMux
    port map (
            O => \N__3222\,
            I => \N__3215\
        );

    \I__563\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3212\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3218\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_12\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3215\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_12\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3212\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_12\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__3205\,
            I => \N__3202\
        );

    \I__558\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3199\,
            I => \N__3194\
        );

    \I__556\ : InMux
    port map (
            O => \N__3198\,
            I => \N__3191\
        );

    \I__555\ : InMux
    port map (
            O => \N__3197\,
            I => \N__3188\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__3194\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_13\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3191\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_13\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3188\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_13\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__3181\,
            I => \N__3177\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__3180\,
            I => \N__3173\
        );

    \I__549\ : InMux
    port map (
            O => \N__3177\,
            I => \N__3170\
        );

    \I__548\ : InMux
    port map (
            O => \N__3176\,
            I => \N__3167\
        );

    \I__547\ : InMux
    port map (
            O => \N__3173\,
            I => \N__3164\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3170\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_14\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3167\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_14\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3164\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_14\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3157\,
            I => \N__3154\
        );

    \I__542\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3151\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3151\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_3_and\
        );

    \I__540\ : InMux
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3145\,
            I => \N__3142\
        );

    \I__538\ : Span4Mux_h
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__537\ : Odrv4
    port map (
            O => \N__3139\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_CO\
        );

    \I__536\ : InMux
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__534\ : Span4Mux_h
    port map (
            O => \N__3130\,
            I => \N__3125\
        );

    \I__533\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3120\
        );

    \I__532\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3120\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__3125\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_15\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3120\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_15\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__528\ : InMux
    port map (
            O => \N__3112\,
            I => \N__3109\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3109\,
            I => \N__3106\
        );

    \I__526\ : Span4Mux_h
    port map (
            O => \N__3106\,
            I => \N__3103\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__3103\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_CO\
        );

    \I__524\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3095\
        );

    \I__523\ : InMux
    port map (
            O => \N__3099\,
            I => \N__3092\
        );

    \I__522\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3089\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3095\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_17\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3092\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_17\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3089\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_17\
        );

    \I__518\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__516\ : Span4Mux_h
    port map (
            O => \N__3076\,
            I => \N__3071\
        );

    \I__515\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3066\
        );

    \I__514\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3066\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__3071\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_16\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3066\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_16\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3061\,
            I => \N__3056\
        );

    \I__510\ : InMux
    port map (
            O => \N__3060\,
            I => \N__3053\
        );

    \I__509\ : InMux
    port map (
            O => \N__3059\,
            I => \N__3050\
        );

    \I__508\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3047\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3053\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_18\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3050\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_18\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3047\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_18\
        );

    \I__504\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3035\
        );

    \I__503\ : InMux
    port map (
            O => \N__3039\,
            I => \N__3032\
        );

    \I__502\ : InMux
    port map (
            O => \N__3038\,
            I => \N__3029\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3035\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_19\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3032\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_19\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3029\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_19\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__3022\,
            I => \N__3019\
        );

    \I__497\ : InMux
    port map (
            O => \N__3019\,
            I => \N__3016\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3016\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_4_and\
        );

    \I__495\ : InMux
    port map (
            O => \N__3013\,
            I => \N__3008\
        );

    \I__494\ : InMux
    port map (
            O => \N__3012\,
            I => \N__3005\
        );

    \I__493\ : InMux
    port map (
            O => \N__3011\,
            I => \N__3002\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3008\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_23\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3005\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_23\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3002\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_23\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__488\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__2989\,
            I => \N__2986\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__2986\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_5_and\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__2983\,
            I => \un1_M_count_q_c2_cascade_\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__2980\,
            I => \un1_M_count_q_c5_cascade_\
        );

    \I__483\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2972\
        );

    \I__482\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2969\
        );

    \I__481\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2966\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2972\,
            I => \N__2961\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2969\,
            I => \N__2961\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__2966\,
            I => \M_count_qZ0Z_6\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__2961\,
            I => \M_count_qZ0Z_6\
        );

    \I__476\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2951\
        );

    \I__475\ : InMux
    port map (
            O => \N__2955\,
            I => \N__2946\
        );

    \I__474\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2946\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__2951\,
            I => \un1_M_count_q_c2\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2946\,
            I => \un1_M_count_q_c2\
        );

    \I__471\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2937\
        );

    \I__470\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2934\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2937\,
            I => \N__2927\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2934\,
            I => \N__2927\
        );

    \I__467\ : InMux
    port map (
            O => \N__2933\,
            I => \N__2922\
        );

    \I__466\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2922\
        );

    \I__465\ : Odrv4
    port map (
            O => \N__2927\,
            I => \M_count_qZ0Z_4\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2922\,
            I => \M_count_qZ0Z_4\
        );

    \I__463\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2914\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2914\,
            I => \un1_M_count_q_c5\
        );

    \I__461\ : InMux
    port map (
            O => \N__2911\,
            I => \N__2905\
        );

    \I__460\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2902\
        );

    \I__459\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2897\
        );

    \I__458\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2897\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2905\,
            I => \N__2894\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2902\,
            I => \N__2891\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2897\,
            I => \M_count_qZ0Z_5\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__2894\,
            I => \M_count_qZ0Z_5\
        );

    \I__453\ : Odrv4
    port map (
            O => \N__2891\,
            I => \M_count_qZ0Z_5\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__2884\,
            I => \N__2881\
        );

    \I__451\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2878\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2878\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_0_and\
        );

    \I__449\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2872\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2872\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_1_and\
        );

    \I__447\ : InMux
    port map (
            O => \N__2869\,
            I => \N__2866\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2866\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_2_and\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__2863\,
            I => \sr_chain_is_sending_0_clk_cascade_\
        );

    \I__444\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2857\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2857\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_1\
        );

    \I__442\ : InMux
    port map (
            O => \N__2854\,
            I => \N__2851\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2851\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_2\
        );

    \I__440\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2845\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_3\
        );

    \I__438\ : InMux
    port map (
            O => \N__2842\,
            I => \N__2838\
        );

    \I__437\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2835\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2838\,
            I => sr_data_to_send_4
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2835\,
            I => sr_data_to_send_4
        );

    \I__434\ : InMux
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2827\,
            I => \N__2824\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__2824\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_4\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__2821\,
            I => \N__2818\
        );

    \I__430\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2814\
        );

    \I__429\ : InMux
    port map (
            O => \N__2817\,
            I => \N__2811\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2814\,
            I => sr_data_to_send_5
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2811\,
            I => sr_data_to_send_5
        );

    \I__426\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2803\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2803\,
            I => \N__2800\
        );

    \I__424\ : Odrv4
    port map (
            O => \N__2800\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_5\
        );

    \I__423\ : InMux
    port map (
            O => \N__2797\,
            I => \N__2793\
        );

    \I__422\ : InMux
    port map (
            O => \N__2796\,
            I => \N__2790\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2793\,
            I => sr_data_to_send_6
        );

    \I__420\ : LocalMux
    port map (
            O => \N__2790\,
            I => sr_data_to_send_6
        );

    \I__419\ : InMux
    port map (
            O => \N__2785\,
            I => \N__2781\
        );

    \I__418\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2778\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2781\,
            I => sr_data_to_send_7
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2778\,
            I => sr_data_to_send_7
        );

    \I__415\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2764\
        );

    \I__414\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2764\
        );

    \I__413\ : InMux
    port map (
            O => \N__2771\,
            I => \N__2761\
        );

    \I__412\ : InMux
    port map (
            O => \N__2770\,
            I => \N__2758\
        );

    \I__411\ : InMux
    port map (
            O => \N__2769\,
            I => \N__2755\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2764\,
            I => \M_count_qZ0Z_0\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2761\,
            I => \M_count_qZ0Z_0\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2758\,
            I => \M_count_qZ0Z_0\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2755\,
            I => \M_count_qZ0Z_0\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__2746\,
            I => \N__2743\
        );

    \I__405\ : InMux
    port map (
            O => \N__2743\,
            I => \N__2740\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2740\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_CO\
        );

    \I__403\ : InMux
    port map (
            O => \N__2737\,
            I => \N__2734\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2734\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_CO\
        );

    \I__401\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2726\
        );

    \I__400\ : InMux
    port map (
            O => \N__2730\,
            I => \N__2723\
        );

    \I__399\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2720\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2726\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_7\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2723\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_7\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2720\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_7\
        );

    \I__395\ : InMux
    port map (
            O => \N__2713\,
            I => \N__2710\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2710\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_CO\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__2707\,
            I => \N__2704\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2704\,
            I => \N__2701\
        );

    \I__391\ : Span4Mux_s1_h
    port map (
            O => \N__2701\,
            I => \N__2698\
        );

    \I__390\ : Sp12to4
    port map (
            O => \N__2698\,
            I => \N__2695\
        );

    \I__389\ : Span12Mux_s11_v
    port map (
            O => \N__2695\,
            I => \N__2692\
        );

    \I__388\ : Span12Mux_h
    port map (
            O => \N__2692\,
            I => \N__2689\
        );

    \I__387\ : Span12Mux_h
    port map (
            O => \N__2689\,
            I => \N__2686\
        );

    \I__386\ : Odrv12
    port map (
            O => \N__2686\,
            I => sr_chain_latch_e1_i
        );

    \I__385\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2680\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2680\,
            I => \un1_M_count_q_axbxc7_m4_0_a2_3\
        );

    \I__383\ : InMux
    port map (
            O => \N__2677\,
            I => \N__2673\
        );

    \I__382\ : InMux
    port map (
            O => \N__2676\,
            I => \N__2670\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2673\,
            I => \M_count_qZ0Z_7\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2670\,
            I => \M_count_qZ0Z_7\
        );

    \I__379\ : InMux
    port map (
            O => \N__2665\,
            I => \N__2662\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2662\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_CO\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__2659\,
            I => \N__2654\
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__2658\,
            I => \N__2651\
        );

    \I__375\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2648\
        );

    \I__374\ : InMux
    port map (
            O => \N__2654\,
            I => \N__2643\
        );

    \I__373\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2643\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2648\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_5\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2643\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_5\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__2638\,
            I => \N__2635\
        );

    \I__369\ : InMux
    port map (
            O => \N__2635\,
            I => \N__2632\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__2629\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_CO\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__2626\,
            I => \N__2623\
        );

    \I__365\ : InMux
    port map (
            O => \N__2623\,
            I => \N__2620\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2620\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_CO\
        );

    \I__363\ : InMux
    port map (
            O => \N__2617\,
            I => \N__2612\
        );

    \I__362\ : InMux
    port map (
            O => \N__2616\,
            I => \N__2609\
        );

    \I__361\ : InMux
    port map (
            O => \N__2615\,
            I => \N__2606\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2612\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_11\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2609\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_11\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2606\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_11\
        );

    \I__357\ : InMux
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2596\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_CO\
        );

    \I__355\ : InMux
    port map (
            O => \N__2593\,
            I => \N__2590\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2590\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_CO\
        );

    \I__353\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2584\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2584\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_CO\
        );

    \I__351\ : InMux
    port map (
            O => \N__2581\,
            I => \N__2578\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2578\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_CO\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__2575\,
            I => \N__2572\
        );

    \I__348\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2569\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2569\,
            I => \N__2566\
        );

    \I__346\ : Odrv4
    port map (
            O => \N__2566\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_CO\
        );

    \I__345\ : InMux
    port map (
            O => \N__2563\,
            I => \N__2558\
        );

    \I__344\ : InMux
    port map (
            O => \N__2562\,
            I => \N__2555\
        );

    \I__343\ : InMux
    port map (
            O => \N__2561\,
            I => \N__2552\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2558\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_6\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2555\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_6\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2552\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_6\
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__2545\,
            I => \N__2542\
        );

    \I__338\ : InMux
    port map (
            O => \N__2542\,
            I => \N__2539\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2539\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_CO\
        );

    \I__336\ : InMux
    port map (
            O => \N__2536\,
            I => \N__2533\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2533\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_CO\
        );

    \I__334\ : InMux
    port map (
            O => \N__2530\,
            I => \N__2525\
        );

    \I__333\ : InMux
    port map (
            O => \N__2529\,
            I => \N__2522\
        );

    \I__332\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2519\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2525\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_1\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2522\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_1\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2519\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_1\
        );

    \I__328\ : InMux
    port map (
            O => \N__2512\,
            I => \N__2509\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2509\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_CO\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2506\,
            I => \N__2501\
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2505\,
            I => \N__2498\
        );

    \I__324\ : InMux
    port map (
            O => \N__2504\,
            I => \N__2495\
        );

    \I__323\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2490\
        );

    \I__322\ : InMux
    port map (
            O => \N__2498\,
            I => \N__2490\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2495\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_2\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2490\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_2\
        );

    \I__319\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2482\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2482\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_CO\
        );

    \I__317\ : InMux
    port map (
            O => \N__2479\,
            I => \N__2474\
        );

    \I__316\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2469\
        );

    \I__315\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2469\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2474\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_3\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2469\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_3\
        );

    \I__312\ : InMux
    port map (
            O => \N__2464\,
            I => \N__2461\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2461\,
            I => \N__2458\
        );

    \I__310\ : Odrv4
    port map (
            O => \N__2458\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_CO\
        );

    \I__309\ : InMux
    port map (
            O => \N__2455\,
            I => \N__2451\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__2454\,
            I => \N__2447\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2451\,
            I => \N__2444\
        );

    \I__306\ : InMux
    port map (
            O => \N__2450\,
            I => \N__2439\
        );

    \I__305\ : InMux
    port map (
            O => \N__2447\,
            I => \N__2439\
        );

    \I__304\ : Odrv4
    port map (
            O => \N__2444\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_10\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2439\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_10\
        );

    \I__302\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2430\
        );

    \I__301\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2426\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2430\,
            I => \N__2423\
        );

    \I__299\ : InMux
    port map (
            O => \N__2429\,
            I => \N__2420\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2426\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_9\
        );

    \I__297\ : Odrv4
    port map (
            O => \N__2423\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_9\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2420\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_9\
        );

    \I__295\ : InMux
    port map (
            O => \N__2413\,
            I => \N__2410\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2410\,
            I => \N__2407\
        );

    \I__293\ : Span4Mux_h
    port map (
            O => \N__2407\,
            I => \N__2404\
        );

    \I__292\ : Odrv4
    port map (
            O => \N__2404\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_CO\
        );

    \I__291\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2398\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2398\,
            I => \N__2393\
        );

    \I__289\ : InMux
    port map (
            O => \N__2397\,
            I => \N__2388\
        );

    \I__288\ : InMux
    port map (
            O => \N__2396\,
            I => \N__2388\
        );

    \I__287\ : Odrv4
    port map (
            O => \N__2393\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_8\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2388\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_8\
        );

    \I__285\ : CascadeMux
    port map (
            O => \N__2383\,
            I => \N__2380\
        );

    \I__284\ : InMux
    port map (
            O => \N__2380\,
            I => \N__2377\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2377\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_CO\
        );

    \I__282\ : InMux
    port map (
            O => \N__2374\,
            I => \N__2369\
        );

    \I__281\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2364\
        );

    \I__280\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2364\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2369\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_4\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2364\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_4\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__2359\,
            I => \N__2341\
        );

    \I__276\ : CascadeMux
    port map (
            O => \N__2358\,
            I => \N__2338\
        );

    \I__275\ : CascadeMux
    port map (
            O => \N__2357\,
            I => \N__2335\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__2356\,
            I => \N__2332\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2355\,
            I => \N__2329\
        );

    \I__272\ : CascadeMux
    port map (
            O => \N__2354\,
            I => \N__2326\
        );

    \I__271\ : CascadeMux
    port map (
            O => \N__2353\,
            I => \N__2323\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__2352\,
            I => \N__2320\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__2351\,
            I => \N__2317\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__2350\,
            I => \N__2314\
        );

    \I__267\ : CascadeMux
    port map (
            O => \N__2349\,
            I => \N__2311\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__2348\,
            I => \N__2308\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__2347\,
            I => \N__2305\
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__2346\,
            I => \N__2302\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__2345\,
            I => \N__2299\
        );

    \I__262\ : CascadeMux
    port map (
            O => \N__2344\,
            I => \N__2296\
        );

    \I__261\ : InMux
    port map (
            O => \N__2341\,
            I => \N__2280\
        );

    \I__260\ : InMux
    port map (
            O => \N__2338\,
            I => \N__2280\
        );

    \I__259\ : InMux
    port map (
            O => \N__2335\,
            I => \N__2280\
        );

    \I__258\ : InMux
    port map (
            O => \N__2332\,
            I => \N__2280\
        );

    \I__257\ : InMux
    port map (
            O => \N__2329\,
            I => \N__2271\
        );

    \I__256\ : InMux
    port map (
            O => \N__2326\,
            I => \N__2271\
        );

    \I__255\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2271\
        );

    \I__254\ : InMux
    port map (
            O => \N__2320\,
            I => \N__2271\
        );

    \I__253\ : InMux
    port map (
            O => \N__2317\,
            I => \N__2262\
        );

    \I__252\ : InMux
    port map (
            O => \N__2314\,
            I => \N__2262\
        );

    \I__251\ : InMux
    port map (
            O => \N__2311\,
            I => \N__2262\
        );

    \I__250\ : InMux
    port map (
            O => \N__2308\,
            I => \N__2262\
        );

    \I__249\ : InMux
    port map (
            O => \N__2305\,
            I => \N__2253\
        );

    \I__248\ : InMux
    port map (
            O => \N__2302\,
            I => \N__2253\
        );

    \I__247\ : InMux
    port map (
            O => \N__2299\,
            I => \N__2253\
        );

    \I__246\ : InMux
    port map (
            O => \N__2296\,
            I => \N__2253\
        );

    \I__245\ : CascadeMux
    port map (
            O => \N__2295\,
            I => \N__2250\
        );

    \I__244\ : CascadeMux
    port map (
            O => \N__2294\,
            I => \N__2247\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2293\,
            I => \N__2244\
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__2292\,
            I => \N__2241\
        );

    \I__241\ : CascadeMux
    port map (
            O => \N__2291\,
            I => \N__2238\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__2290\,
            I => \N__2235\
        );

    \I__239\ : CascadeMux
    port map (
            O => \N__2289\,
            I => \N__2232\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2280\,
            I => \N__2227\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2271\,
            I => \N__2227\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2262\,
            I => \N__2222\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2253\,
            I => \N__2222\
        );

    \I__234\ : InMux
    port map (
            O => \N__2250\,
            I => \N__2215\
        );

    \I__233\ : InMux
    port map (
            O => \N__2247\,
            I => \N__2215\
        );

    \I__232\ : InMux
    port map (
            O => \N__2244\,
            I => \N__2215\
        );

    \I__231\ : InMux
    port map (
            O => \N__2241\,
            I => \N__2206\
        );

    \I__230\ : InMux
    port map (
            O => \N__2238\,
            I => \N__2206\
        );

    \I__229\ : InMux
    port map (
            O => \N__2235\,
            I => \N__2206\
        );

    \I__228\ : InMux
    port map (
            O => \N__2232\,
            I => \N__2206\
        );

    \I__227\ : Odrv12
    port map (
            O => \N__2227\,
            I => \CONSTANT_ONE_NET\
        );

    \I__226\ : Odrv4
    port map (
            O => \N__2222\,
            I => \CONSTANT_ONE_NET\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2215\,
            I => \CONSTANT_ONE_NET\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2206\,
            I => \CONSTANT_ONE_NET\
        );

    \I__223\ : InMux
    port map (
            O => \N__2197\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1\
        );

    \I__222\ : InMux
    port map (
            O => \N__2194\,
            I => \bfn_26_21_0_\
        );

    \I__221\ : CascadeMux
    port map (
            O => \N__2191\,
            I => \un1_M_count_q_axbxc7_m4_0_a2_2_cascade_\
        );

    \I__220\ : InMux
    port map (
            O => \N__2188\,
            I => \N__2185\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__2185\,
            I => \N__2182\
        );

    \I__218\ : Odrv4
    port map (
            O => \N__2182\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_CO\
        );

    \I__217\ : InMux
    port map (
            O => \N__2179\,
            I => \N__2175\
        );

    \I__216\ : InMux
    port map (
            O => \N__2178\,
            I => \N__2172\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__2175\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_0\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__2172\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_0\
        );

    \I__213\ : InMux
    port map (
            O => \N__2167\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1\
        );

    \I__212\ : InMux
    port map (
            O => \N__2164\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1\
        );

    \I__211\ : InMux
    port map (
            O => \N__2161\,
            I => \bfn_26_20_0_\
        );

    \I__210\ : InMux
    port map (
            O => \N__2158\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1\
        );

    \I__209\ : InMux
    port map (
            O => \N__2155\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1\
        );

    \I__208\ : InMux
    port map (
            O => \N__2152\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1\
        );

    \I__207\ : InMux
    port map (
            O => \N__2149\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1\
        );

    \I__206\ : InMux
    port map (
            O => \N__2146\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1\
        );

    \I__205\ : InMux
    port map (
            O => \N__2143\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1\
        );

    \I__204\ : InMux
    port map (
            O => \N__2140\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1\
        );

    \I__203\ : InMux
    port map (
            O => \N__2137\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1\
        );

    \I__202\ : InMux
    port map (
            O => \N__2134\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1\
        );

    \I__201\ : InMux
    port map (
            O => \N__2131\,
            I => \bfn_26_19_0_\
        );

    \I__200\ : InMux
    port map (
            O => \N__2128\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1\
        );

    \I__199\ : InMux
    port map (
            O => \N__2125\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1\
        );

    \I__198\ : InMux
    port map (
            O => \N__2122\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1\
        );

    \I__197\ : InMux
    port map (
            O => \N__2119\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1\
        );

    \I__196\ : InMux
    port map (
            O => \N__2116\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1\
        );

    \I__195\ : InMux
    port map (
            O => \N__2113\,
            I => \N__2110\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__2110\,
            I => \reset_cond.M_stage_qZ0Z_1\
        );

    \I__193\ : InMux
    port map (
            O => \N__2107\,
            I => \N__2104\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__2104\,
            I => \reset_cond.M_stage_qZ0Z_0\
        );

    \I__191\ : InMux
    port map (
            O => \N__2101\,
            I => \N__2089\
        );

    \I__190\ : InMux
    port map (
            O => \N__2100\,
            I => \N__2089\
        );

    \I__189\ : InMux
    port map (
            O => \N__2099\,
            I => \N__2089\
        );

    \I__188\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2089\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__2089\,
            I => \N__2086\
        );

    \I__186\ : Span12Mux_v
    port map (
            O => \N__2086\,
            I => \N__2083\
        );

    \I__185\ : Odrv12
    port map (
            O => \N__2083\,
            I => rst_n_c
        );

    \I__184\ : InMux
    port map (
            O => \N__2080\,
            I => \N__2077\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__2077\,
            I => \reset_cond.M_stage_qZ0Z_2\
        );

    \I__182\ : InMux
    port map (
            O => \N__2074\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1\
        );

    \I__181\ : InMux
    port map (
            O => \N__2071\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1\
        );

    \I__180\ : InMux
    port map (
            O => \N__2068\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1\
        );

    \I__179\ : InMux
    port map (
            O => \N__2065\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1\
        );

    \IN_MUX_bfv_28_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_28_17_0_\
        );

    \IN_MUX_bfv_29_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_29_18_0_\
        );

    \IN_MUX_bfv_26_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_26_18_0_\
        );

    \IN_MUX_bfv_26_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1\,
            carryinitout => \bfn_26_19_0_\
        );

    \IN_MUX_bfv_26_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1\,
            carryinitout => \bfn_26_20_0_\
        );

    \IN_MUX_bfv_26_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1\,
            carryinitout => \bfn_26_21_0_\
        );

    \IN_MUX_bfv_30_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_30_15_0_\
        );

    \IN_MUX_bfv_30_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_main_clock_count_q_1_cry_7\,
            carryinitout => \bfn_30_16_0_\
        );

    \IN_MUX_bfv_30_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_main_clock_count_q_1_cry_15\,
            carryinitout => \bfn_30_17_0_\
        );

    \IN_MUX_bfv_30_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_main_clock_count_q_1_cry_23\,
            carryinitout => \bfn_30_18_0_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3700\,
            GLOBALBUFFEROUTPUT => \sr_chain.N_44_g\
        );

    \reset_cond.M_stage_q_RNIFG9D_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4696\,
            GLOBALBUFFEROUTPUT => \N_108_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \reset_cond.M_stage_q_1_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2107\,
            lcout => \reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_2_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2100\,
            in2 => \_gnd_net_\,
            in3 => \N__2113\,
            lcout => \reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_0_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_3_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2101\,
            in2 => \_gnd_net_\,
            in3 => \N__2080\,
            lcout => \M_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_26_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_0_LC_26_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__4949\,
            in1 => \N__2179\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_26_18_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1\,
            clk => \N__4750\,
            ce => 'H',
            sr => \N__3454\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_LUT4_0_LC_26_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2529\,
            in2 => \N__2289\,
            in3 => \N__2074\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_0_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_LUT4_0_LC_26_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2504\,
            in2 => \N__2293\,
            in3 => \N__2071\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_1_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_LUT4_0_LC_26_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2479\,
            in2 => \N__2290\,
            in3 => \N__2068\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_2_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_LUT4_0_LC_26_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2374\,
            in2 => \N__2294\,
            in3 => \N__2065\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_3_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_LUT4_0_LC_26_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2657\,
            in2 => \N__2291\,
            in3 => \N__2140\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_4_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_LUT4_0_LC_26_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2562\,
            in2 => \N__2295\,
            in3 => \N__2137\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_5_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_LUT4_0_LC_26_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2730\,
            in2 => \N__2292\,
            in3 => \N__2134\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_6_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_LUT4_0_LC_26_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2401\,
            in2 => \N__2350\,
            in3 => \N__2131\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_7_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_26_19_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_LUT4_0_LC_26_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2434\,
            in2 => \N__2347\,
            in3 => \N__2128\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_8_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_LUT4_0_LC_26_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2455\,
            in2 => \N__2351\,
            in3 => \N__2125\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_9_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_LUT4_0_LC_26_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2616\,
            in2 => \N__2344\,
            in3 => \N__2122\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_10_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_LUT4_0_LC_26_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3222\,
            in2 => \N__2348\,
            in3 => \N__2119\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_11_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_LUT4_0_LC_26_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3198\,
            in2 => \N__2345\,
            in3 => \N__2116\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_12_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_LUT4_0_LC_26_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3176\,
            in2 => \N__2349\,
            in3 => \N__2167\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_13_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_LUT4_0_LC_26_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3136\,
            in2 => \N__2346\,
            in3 => \N__2164\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_14_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_LUT4_0_LC_26_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3082\,
            in2 => \N__2352\,
            in3 => \N__2161\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_15_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_26_20_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_LUT4_0_LC_26_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3099\,
            in2 => \N__2356\,
            in3 => \N__2158\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_16_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_LUT4_0_LC_26_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3059\,
            in2 => \N__2353\,
            in3 => \N__2155\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_17_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_LUT4_0_LC_26_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3039\,
            in2 => \N__2357\,
            in3 => \N__2152\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_18_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_LUT4_0_LC_26_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3517\,
            in2 => \N__2354\,
            in3 => \N__2149\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_19_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_LUT4_0_LC_26_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3481\,
            in2 => \N__2358\,
            in3 => \N__2146\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_20_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_LUT4_0_LC_26_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3550\,
            in2 => \N__2355\,
            in3 => \N__2143\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_21_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_LUT4_0_LC_26_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3012\,
            in2 => \N__2359\,
            in3 => \N__2197\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_22_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_LUT4_0_LC_26_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2194\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_11_cry_23_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNO_1_7_LC_27_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3368\,
            in1 => \N__3421\,
            in2 => \N__3324\,
            in3 => \N__2770\,
            lcout => OPEN,
            ltout => \un1_M_count_q_axbxc7_m4_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNO_0_7_LC_27_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2977\,
            in1 => \N__2911\,
            in2 => \N__2191\,
            in3 => \N__2941\,
            lcout => \un1_M_count_q_axbxc7_m4_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_1_LC_27_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__4951\,
            in1 => \N__3425\,
            in2 => \N__4531\,
            in3 => \N__2773\,
            lcout => \M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4746\,
            ce => 'H',
            sr => \N__4694\
        );

    \M_count_q_3_LC_27_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__2955\,
            in1 => \_gnd_net_\,
            in2 => \N__3380\,
            in3 => \N__3320\,
            lcout => \M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4746\,
            ce => 'H',
            sr => \N__4694\
        );

    \M_count_q_2_LC_27_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3370\,
            in2 => \_gnd_net_\,
            in3 => \N__2954\,
            lcout => \M_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4746\,
            ce => 'H',
            sr => \N__4694\
        );

    \M_count_q_0_LC_27_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__2772\,
            in1 => \N__4524\,
            in2 => \_gnd_net_\,
            in3 => \N__4952\,
            lcout => \M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4746\,
            ce => 'H',
            sr => \N__4694\
        );

    \sr_chain.M_sr_rest_cycles_q_9_LC_27_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__2188\,
            in1 => \N__3628\,
            in2 => \_gnd_net_\,
            in3 => \N__2433\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4748\,
            ce => 'H',
            sr => \N__3460\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_RNO_LC_27_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2528\,
            in1 => \N__2178\,
            in2 => \N__2505\,
            in3 => \N__2477\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_1_LC_27_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__2530\,
            in1 => \N__2536\,
            in2 => \_gnd_net_\,
            in3 => \N__3617\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4751\,
            ce => 'H',
            sr => \N__3458\
        );

    \sr_chain.M_sr_rest_cycles_q_2_LC_27_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001011010010"
        )
    port map (
            in0 => \N__3618\,
            in1 => \N__2512\,
            in2 => \N__2506\,
            in3 => \_gnd_net_\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4751\,
            ce => 'H',
            sr => \N__3458\
        );

    \sr_chain.M_sr_rest_cycles_q_3_LC_27_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__2478\,
            in1 => \N__2485\,
            in2 => \_gnd_net_\,
            in3 => \N__3619\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4751\,
            ce => 'H',
            sr => \N__3458\
        );

    \sr_chain.M_sr_rest_cycles_q_10_LC_27_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2450\,
            in2 => \N__3626\,
            in3 => \N__2464\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4751\,
            ce => 'H',
            sr => \N__3458\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_RNO_LC_27_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2396\,
            in1 => \N__2615\,
            in2 => \N__2454\,
            in3 => \N__2429\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_8_LC_27_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2397\,
            in2 => \N__3627\,
            in3 => \N__2413\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4751\,
            ce => 'H',
            sr => \N__3458\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_RNO_LC_27_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2561\,
            in1 => \N__2729\,
            in2 => \N__2658\,
            in3 => \N__2372\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_4_LC_27_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010110101010"
        )
    port map (
            in0 => \N__2373\,
            in1 => \_gnd_net_\,
            in2 => \N__2383\,
            in3 => \N__3598\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4755\,
            ce => 'H',
            sr => \N__3457\
        );

    \sr_chain.M_sr_rest_cycles_q_5_LC_27_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001011010010"
        )
    port map (
            in0 => \N__3599\,
            in1 => \N__2665\,
            in2 => \N__2659\,
            in3 => \_gnd_net_\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4755\,
            ce => 'H',
            sr => \N__3457\
        );

    \sr_chain.M_sr_rest_cycles_q_24_LC_27_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010001101"
        )
    port map (
            in0 => \N__4940\,
            in1 => \N__4122\,
            in2 => \N__2638\,
            in3 => \N__3250\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4755\,
            ce => 'H',
            sr => \N__3457\
        );

    \sr_chain.M_sr_rest_cycles_q_11_LC_27_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__4120\,
            in1 => \N__2617\,
            in2 => \N__2626\,
            in3 => \N__4941\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4755\,
            ce => 'H',
            sr => \N__3457\
        );

    \sr_chain.M_sr_rest_cycles_q_12_LC_27_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010101101"
        )
    port map (
            in0 => \N__4939\,
            in1 => \N__4121\,
            in2 => \N__3226\,
            in3 => \N__2599\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4755\,
            ce => 'H',
            sr => \N__3457\
        );

    \sr_chain.M_sr_rest_cycles_q_13_LC_27_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011000011"
        )
    port map (
            in0 => \N__4105\,
            in1 => \N__2593\,
            in2 => \N__3205\,
            in3 => \N__4936\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4758\,
            ce => 'H',
            sr => \N__3455\
        );

    \sr_chain.M_sr_rest_cycles_q_14_LC_27_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010101101"
        )
    port map (
            in0 => \N__4934\,
            in1 => \N__4106\,
            in2 => \N__3181\,
            in3 => \N__2587\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4758\,
            ce => 'H',
            sr => \N__3455\
        );

    \sr_chain.M_sr_rest_cycles_q_17_LC_27_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__2581\,
            in1 => \N__3595\,
            in2 => \_gnd_net_\,
            in3 => \N__3100\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4758\,
            ce => 'H',
            sr => \N__3455\
        );

    \sr_chain.M_sr_rest_cycles_q_6_LC_27_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__4109\,
            in1 => \N__2563\,
            in2 => \N__2575\,
            in3 => \N__4938\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4758\,
            ce => 'H',
            sr => \N__3455\
        );

    \sr_chain.M_sr_rest_cycles_q_19_LC_27_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010001101"
        )
    port map (
            in0 => \N__4935\,
            in1 => \N__4108\,
            in2 => \N__2545\,
            in3 => \N__3040\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4758\,
            ce => 'H',
            sr => \N__3455\
        );

    \sr_chain.M_sr_rest_cycles_q_18_LC_27_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__4107\,
            in1 => \N__3060\,
            in2 => \N__2746\,
            in3 => \N__4937\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4758\,
            ce => 'H',
            sr => \N__3455\
        );

    \sr_chain.M_sr_rest_cycles_q_7_LC_27_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__2737\,
            in1 => \N__3596\,
            in2 => \_gnd_net_\,
            in3 => \N__2731\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4758\,
            ce => 'H',
            sr => \N__3455\
        );

    \sr_chain.M_sr_rest_cycles_q_23_LC_27_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__2713\,
            in1 => \N__3597\,
            in2 => \_gnd_net_\,
            in3 => \N__3013\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4761\,
            ce => 'H',
            sr => \N__3453\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIH9O82_LC_27_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4950\,
            in2 => \_gnd_net_\,
            in3 => \N__4123\,
            lcout => sr_chain_latch_e1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_7_LC_28_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__4932\,
            in1 => \N__2677\,
            in2 => \N__4510\,
            in3 => \N__2683\,
            lcout => \M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4747\,
            ce => 'H',
            sr => \N__4695\
        );

    \M_count_q_RNIR63U_7_LC_28_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2785\,
            in1 => \N__2676\,
            in2 => \_gnd_net_\,
            in3 => \N__3286\,
            lcout => sr_data_to_send_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIQ53U_6_LC_28_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__3285\,
            in1 => \N__2976\,
            in2 => \_gnd_net_\,
            in3 => \N__2797\,
            lcout => sr_data_to_send_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIO33U_4_LC_28_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2940\,
            in1 => \N__3283\,
            in2 => \_gnd_net_\,
            in3 => \N__2842\,
            lcout => sr_data_to_send_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIP43U_5_LC_28_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__3284\,
            in1 => \N__2910\,
            in2 => \N__2821\,
            in3 => \_gnd_net_\,
            lcout => sr_data_to_send_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_is_sending_q_RNI73BG_0_LC_28_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4493\,
            in2 => \_gnd_net_\,
            in3 => \N__4931\,
            lcout => sr_chain_is_sending_0_clk,
            ltout => \sr_chain_is_sending_0_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIKV2U_0_LC_28_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2771\,
            in2 => \N__2863\,
            in3 => \N__3657\,
            lcout => sr_data_to_send_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_data_buffer_q_esr_1_LC_28_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3639\,
            in1 => \N__3396\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4749\,
            ce => \N__3670\,
            sr => \N__4693\
        );

    \sr_chain.M_sr_data_buffer_q_esr_2_LC_28_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3336\,
            in1 => \N__2860\,
            in2 => \_gnd_net_\,
            in3 => \N__4530\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4749\,
            ce => \N__3670\,
            sr => \N__4693\
        );

    \sr_chain.M_sr_data_buffer_q_esr_3_LC_28_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3261\,
            in1 => \N__2854\,
            in2 => \_gnd_net_\,
            in3 => \N__4485\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4749\,
            ce => \N__3670\,
            sr => \N__4693\
        );

    \sr_chain.M_sr_data_buffer_q_esr_4_LC_28_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2848\,
            in1 => \N__4528\,
            in2 => \_gnd_net_\,
            in3 => \N__2841\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4749\,
            ce => \N__3670\,
            sr => \N__4693\
        );

    \sr_chain.M_sr_data_buffer_q_esr_5_LC_28_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2830\,
            in1 => \N__4482\,
            in2 => \_gnd_net_\,
            in3 => \N__2817\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4749\,
            ce => \N__3670\,
            sr => \N__4693\
        );

    \sr_chain.M_sr_data_buffer_q_esr_6_LC_28_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2806\,
            in1 => \N__4529\,
            in2 => \_gnd_net_\,
            in3 => \N__2796\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4749\,
            ce => \N__3670\,
            sr => \N__4693\
        );

    \sr_chain.M_sr_data_buffer_q_esr_7_LC_28_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4587\,
            in1 => \N__4483\,
            in2 => \_gnd_net_\,
            in3 => \N__2784\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4749\,
            ce => \N__3670\,
            sr => \N__4693\
        );

    \M_count_q_RNI2TQB1_1_LC_28_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2769\,
            in1 => \N__4479\,
            in2 => \N__3426\,
            in3 => \N__4881\,
            lcout => \un1_M_count_q_c2\,
            ltout => \un1_M_count_q_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIIR2L2_4_LC_28_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2932\,
            in1 => \N__3318\,
            in2 => \N__2983\,
            in3 => \N__3369\,
            lcout => \un1_M_count_q_c5\,
            ltout => \un1_M_count_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_6_LC_28_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2909\,
            in2 => \N__2980\,
            in3 => \N__2975\,
            lcout => \M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4752\,
            ce => 'H',
            sr => \N__4692\
        );

    \M_count_q_4_LC_28_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__2933\,
            in1 => \N__3319\,
            in2 => \N__3385\,
            in3 => \N__2956\,
            lcout => \M_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4752\,
            ce => 'H',
            sr => \N__4692\
        );

    \M_count_q_5_LC_28_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2908\,
            in2 => \_gnd_net_\,
            in3 => \N__2917\,
            lcout => \M_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4752\,
            ce => 'H',
            sr => \N__4692\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_LC_28_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2884\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_28_17_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_LC_28_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2875\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_0\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_LC_28_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2869\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_LC_28_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3157\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_2\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_LC_28_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3022\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_3\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_LC_28_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2995\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_4\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_inv_LC_28_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3238\,
            in3 => \N__3249\,
            lcout => \sr_chain.M_sr_rest_cycles_q_i_24\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_5\,
            carryout => \sr_chain_un1_M_sr_rest_cycles_q_1_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_LUT4_0_LC_28_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3229\,
            lcout => \sr_chain_un1_M_sr_rest_cycles_q_1_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_RNO_LC_28_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3221\,
            in1 => \N__3197\,
            in2 => \N__3180\,
            in3 => \N__3128\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_15_LC_28_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__3129\,
            in1 => \N__3148\,
            in2 => \_gnd_net_\,
            in3 => \N__3594\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4759\,
            ce => 'H',
            sr => \N__3459\
        );

    \sr_chain.M_sr_rest_cycles_q_16_LC_28_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010100101"
        )
    port map (
            in0 => \N__3075\,
            in1 => \N__4101\,
            in2 => \N__3115\,
            in3 => \N__4907\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4759\,
            ce => 'H',
            sr => \N__3459\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_RNO_LC_28_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3098\,
            in1 => \N__3074\,
            in2 => \N__3061\,
            in3 => \N__3038\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_RNO_LC_28_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3545\,
            in1 => \N__3476\,
            in2 => \N__3516\,
            in3 => \N__3011\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIFAS5_LC_28_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4933\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_22_LC_28_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__4104\,
            in1 => \N__3549\,
            in2 => \N__3562\,
            in3 => \N__4944\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4763\,
            ce => 'H',
            sr => \N__3456\
        );

    \sr_chain.M_sr_rest_cycles_q_20_LC_28_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__4102\,
            in1 => \N__3515\,
            in2 => \N__3529\,
            in3 => \N__4942\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4763\,
            ce => 'H',
            sr => \N__3456\
        );

    \sr_chain.M_sr_rest_cycles_q_21_LC_28_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__4103\,
            in1 => \N__3480\,
            in2 => \N__3493\,
            in3 => \N__4943\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4763\,
            ce => 'H',
            sr => \N__3456\
        );

    \M_count_q_RNIL03U_1_LC_29_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3397\,
            in1 => \N__3430\,
            in2 => \_gnd_net_\,
            in3 => \N__3287\,
            lcout => sr_data_to_send_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIM13U_2_LC_29_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__3288\,
            in1 => \N__3384\,
            in2 => \_gnd_net_\,
            in3 => \N__3337\,
            lcout => sr_data_to_send_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIN23U_3_LC_29_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3325\,
            in1 => \N__3289\,
            in2 => \_gnd_net_\,
            in3 => \N__3262\,
            lcout => sr_data_to_send_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_4_c_RNO_LC_29_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4236\,
            in1 => \N__4200\,
            in2 => \N__4258\,
            in3 => \N__4185\,
            lcout => \sr_chain.M_main_clock_count_d8_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_RNIL1D81_1_LC_29_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4008\,
            in1 => \_gnd_net_\,
            in2 => \N__3688\,
            in3 => \N__3716\,
            lcout => \sr_chain.un1_M_sr_clock_count_q_1_c2\,
            ltout => \sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_2_LC_29_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__3884\,
            in1 => \_gnd_net_\,
            in2 => \N__3691\,
            in3 => \N__3932\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_3_c_RNO_LC_29_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3847\,
            in1 => \N__4272\,
            in2 => \N__3832\,
            in3 => \N__3813\,
            lcout => \sr_chain.M_main_clock_count_d8_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_1_LC_29_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__3718\,
            in1 => \N__3687\,
            in2 => \N__3888\,
            in3 => \N__4010\,
            lcout => \sr_chain.M_sr_clock_count_qZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_RNI74IL_3_LC_29_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3902\,
            lcout => OPEN,
            ltout => \sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_RNIV7TL1_1_LC_29_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__3950\,
            in1 => \N__3683\,
            in2 => \N__3673\,
            in3 => \N__4007\,
            lcout => \sr_chain.un1_M_sr_clock_count_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_0_LC_29_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4009\,
            in1 => \N__3880\,
            in2 => \_gnd_net_\,
            in3 => \N__3717\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNIIHTA1_LC_29_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__4662\,
            in1 => \N__3726\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_data_buffer_q_0_LC_29_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__4480\,
            in1 => \N__3727\,
            in2 => \N__3643\,
            in3 => \N__3658\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4756\,
            ce => 'H',
            sr => \N__4684\
        );

    \sr_chain.M_sr_is_sending_q_LC_29_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110011011101110"
        )
    port map (
            in0 => \N__4854\,
            in1 => \N__4481\,
            in2 => \N__4573\,
            in3 => \N__4060\,
            lcout => sr_chain_latch13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4756\,
            ce => 'H',
            sr => \N__4684\
        );

    \sr_chain.M_sr_is_sending_q_RNI73BG_LC_29_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4454\,
            in2 => \_gnd_net_\,
            in3 => \N__4853\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNI31KT_LC_29_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010100000000"
        )
    port map (
            in0 => \N__4486\,
            in1 => \N__4059\,
            in2 => \N__4027\,
            in3 => \N__4914\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_1_c_RNO_LC_29_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4332\,
            in1 => \N__4302\,
            in2 => \N__4366\,
            in3 => \N__4287\,
            lcout => \sr_chain.M_main_clock_count_d8_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_is_sending_q_RNIMJKT_LC_29_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__4661\,
            in1 => \_gnd_net_\,
            in2 => \N__4509\,
            in3 => \N__4916\,
            lcout => \sr_chain.M_sr_is_sending_q_RNIMJKTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_0_c_RNO_LC_29_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4380\,
            in1 => \N__4137\,
            in2 => \N__4222\,
            in3 => \N__4395\,
            lcout => \sr_chain.M_main_clock_count_d8_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNII1RI_LC_29_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4915\,
            in2 => \N__4508\,
            in3 => \N__4058\,
            lcout => \sr_chain.M_main_clock_count_d_0_sqmuxa\,
            ltout => \sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_LC_29_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3703\,
            in3 => \N__4660\,
            lcout => \sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_5_c_RNO_LC_29_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4317\,
            in1 => \N__4347\,
            in2 => \N__4171\,
            in3 => \N__4152\,
            lcout => \sr_chain.M_main_clock_count_d8_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_2_c_RNO_LC_29_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5059\,
            in1 => \N__4989\,
            in2 => \N__5026\,
            in3 => \N__5040\,
            lcout => \sr_chain.M_main_clock_count_d8_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_0_c_LC_29_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3799\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_29_18_0_\,
            carryout => \sr_chain.M_main_clock_count_d8_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_1_c_LC_29_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3790\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_0\,
            carryout => \sr_chain.M_main_clock_count_d8_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_2_c_LC_29_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3781\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_1\,
            carryout => \sr_chain.M_main_clock_count_d8_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_3_c_LC_29_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_2\,
            carryout => \sr_chain.M_main_clock_count_d8_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_4_c_LC_29_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3760\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_3\,
            carryout => \sr_chain.M_main_clock_count_d8_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_5_c_LC_29_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_4\,
            carryout => \sr_chain.M_main_clock_count_d8_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_inv_LC_29_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3739\,
            in3 => \N__5007\,
            lcout => \sr_chain.M_main_clock_count_q_i_23\,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_5\,
            carryout => \sr_chain.M_main_clock_count_d8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_THRU_LUT4_0_LC_29_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3730\,
            lcout => \sr_chain.M_main_clock_count_d8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_bit_q_RNO_0_LC_29_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__4022\,
            in1 => \N__4498\,
            in2 => \N__3964\,
            in3 => \N__4053\,
            lcout => \sr_chain.M_sr_bit_d_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNI2VR22_LC_29_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__4570\,
            in1 => \N__4497\,
            in2 => \_gnd_net_\,
            in3 => \N__4052\,
            lcout => \sr_chain.latch_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNIPG9U1_LC_29_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__4054\,
            in1 => \N__4571\,
            in2 => \_gnd_net_\,
            in3 => \N__4945\,
            lcout => OPEN,
            ltout => \sr_chain.M_sr_bit_d12_m_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_RNIHJDP2_0_LC_29_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100110011"
        )
    port map (
            in0 => \N__4023\,
            in1 => \N__4954\,
            in2 => \N__3985\,
            in3 => \N__4499\,
            lcout => sr_clk_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_4_LC_30_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__3913\,
            in1 => \N__3904\,
            in2 => \N__3960\,
            in3 => \N__3934\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4754\,
            ce => 'H',
            sr => \N__3889\
        );

    \sr_chain.M_sr_clock_count_q_3_LC_30_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__3903\,
            in1 => \N__3933\,
            in2 => \_gnd_net_\,
            in3 => \N__3912\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4754\,
            ce => 'H',
            sr => \N__3889\
        );

    \sr_chain.M_main_clock_count_q_0_LC_30_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3846\,
            in2 => \N__3862\,
            in3 => \N__3861\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_30_15_0_\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_0\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_1_LC_30_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3831\,
            in2 => \_gnd_net_\,
            in3 => \N__3817\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_0\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_1\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_2_LC_30_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3814\,
            in2 => \_gnd_net_\,
            in3 => \N__3802\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_1\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_2\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_3_LC_30_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4273\,
            in2 => \_gnd_net_\,
            in3 => \N__4261\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_2\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_3\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_4_LC_30_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4254\,
            in2 => \_gnd_net_\,
            in3 => \N__4240\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_3\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_4\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_5_LC_30_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4237\,
            in2 => \_gnd_net_\,
            in3 => \N__4225\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_4\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_5\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_6_LC_30_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4218\,
            in2 => \_gnd_net_\,
            in3 => \N__4204\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_5\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_6\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_7_LC_30_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4201\,
            in2 => \_gnd_net_\,
            in3 => \N__4189\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_6\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_7\,
            clk => \N__4757\,
            ce => 'H',
            sr => \N__4978\
        );

    \sr_chain.M_main_clock_count_q_8_LC_30_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4186\,
            in2 => \_gnd_net_\,
            in3 => \N__4174\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_30_16_0_\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_8\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_9_LC_30_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4170\,
            in2 => \_gnd_net_\,
            in3 => \N__4156\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_8\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_9\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_10_LC_30_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4153\,
            in2 => \_gnd_net_\,
            in3 => \N__4141\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_9\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_10\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_11_LC_30_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4138\,
            in2 => \_gnd_net_\,
            in3 => \N__4126\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_10\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_11\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_12_LC_30_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4396\,
            in2 => \_gnd_net_\,
            in3 => \N__4384\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_11\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_12\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_13_LC_30_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4381\,
            in2 => \_gnd_net_\,
            in3 => \N__4369\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_12\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_13\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_14_LC_30_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4365\,
            in2 => \_gnd_net_\,
            in3 => \N__4351\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_14\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_13\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_14\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_15_LC_30_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4348\,
            in2 => \_gnd_net_\,
            in3 => \N__4336\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_15\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_14\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_15\,
            clk => \N__4760\,
            ce => 'H',
            sr => \N__4976\
        );

    \sr_chain.M_main_clock_count_q_16_LC_30_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4333\,
            in2 => \_gnd_net_\,
            in3 => \N__4321\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_30_17_0_\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_16\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_17_LC_30_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4318\,
            in2 => \_gnd_net_\,
            in3 => \N__4306\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_17\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_16\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_17\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_18_LC_30_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4303\,
            in2 => \_gnd_net_\,
            in3 => \N__4291\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_18\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_17\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_18\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_19_LC_30_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4288\,
            in2 => \_gnd_net_\,
            in3 => \N__4276\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_19\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_18\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_19\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_20_LC_30_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5058\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_20\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_19\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_20\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_21_LC_30_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5041\,
            in2 => \_gnd_net_\,
            in3 => \N__5029\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_21\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_20\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_21\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_22_LC_30_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5025\,
            in2 => \_gnd_net_\,
            in3 => \N__5011\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_22\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_21\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_22\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_23_LC_30_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5008\,
            in2 => \_gnd_net_\,
            in3 => \N__4996\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_23\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_22\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_23\,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4975\
        );

    \sr_chain.M_main_clock_count_q_24_LC_30_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4990\,
            in2 => \_gnd_net_\,
            in3 => \N__4993\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4764\,
            ce => 'H',
            sr => \N__4977\
        );

    \sr_chain.M_sr_bit_q_LC_30_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__4408\,
            in1 => \N__4960\,
            in2 => \N__4782\,
            in3 => \N__4953\,
            lcout => sr_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4765\,
            ce => 'H',
            sr => \N__4688\
        );

    \sr_chain.M_sr_bit_q_RNO_1_LC_31_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__4588\,
            in1 => \N__4572\,
            in2 => \N__4543\,
            in3 => \N__4511\,
            lcout => \sr_chain.M_sr_bit_q_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
