-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Oct 23 2022 18:16:08

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    led : out std_logic_vector(7 downto 0);
    usb_tx : out std_logic;
    trigger : in std_logic;
    rst_n : in std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2047\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2029\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2008\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1941\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1935\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1921\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1893\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1865\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1834\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1810\ : std_logic;
signal \N__1807\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1803\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1801\ : std_logic;
signal \N__1800\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1796\ : std_logic;
signal \N__1785\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1777\ : std_logic;
signal \N__1774\ : std_logic;
signal \N__1771\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1764\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1738\ : std_logic;
signal \N__1735\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1722\ : std_logic;
signal \N__1719\ : std_logic;
signal \N__1716\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1708\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1704\ : std_logic;
signal \N__1701\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1674\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1666\ : std_logic;
signal \N__1663\ : std_logic;
signal \N__1660\ : std_logic;
signal \N__1657\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1650\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1641\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1630\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1591\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1586\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1575\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1567\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1558\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1546\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1525\ : std_logic;
signal \N__1524\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1521\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1498\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1483\ : std_logic;
signal \N__1480\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1470\ : std_logic;
signal \N__1467\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1450\ : std_logic;
signal \N__1447\ : std_logic;
signal \N__1444\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1438\ : std_logic;
signal \N__1435\ : std_logic;
signal \N__1432\ : std_logic;
signal \N__1429\ : std_logic;
signal \N__1426\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1423\ : std_logic;
signal \N__1414\ : std_logic;
signal \N__1411\ : std_logic;
signal \N__1408\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1404\ : std_logic;
signal \N__1401\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1393\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \un1_M_count_q_ac0_1_cascade_\ : std_logic;
signal \un1_M_count_q_ac0_1\ : std_logic;
signal \click_dtct_out3_cascade_\ : std_logic;
signal \un1_M_count_q_ac0_7_cascade_\ : std_logic;
signal click_dtct_out_d : std_logic;
signal \click_dtct_out_d_cascade_\ : std_logic;
signal \un1_M_count_q_ac0_7\ : std_logic;
signal \uart_tx.N_134_i_cascade_\ : std_logic;
signal \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\ : std_logic;
signal \uart_tx.N_182_0_cascade_\ : std_logic;
signal \uart_tx.N_143_0_cascade_\ : std_logic;
signal \uart_tx_N_185_cascade_\ : std_logic;
signal \click_dtct_M_count_d6_0_1_cascade_\ : std_logic;
signal \uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_\ : std_logic;
signal \uart_tx_N_187\ : std_logic;
signal \un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_\ : std_logic;
signal \un1_M_count_q_ac0_5_m2_0_a2_3\ : std_logic;
signal \un1_M_count_q_ac0_5_m2_0_a2_3_cascade_\ : std_logic;
signal \un1_M_count_q_ac0_out\ : std_logic;
signal click_dtct_out3 : std_logic;
signal \M_reset_cond_out_0\ : std_logic;
signal \un1_M_count_q_axbxc7_1\ : std_logic;
signal \btn_cond.out_17_6_cascade_\ : std_logic;
signal \btn_cond.out_17_8\ : std_logic;
signal \btn_cond_out_17_cascade_\ : std_logic;
signal click_dtct_out8 : std_logic;
signal \btn_cond.out_17_7\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal rst_n_c : std_logic;
signal \reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \uart_tx.N_186_1_i\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_0\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \uart_tx.M_ctr_qZ1Z_1\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_0\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_2\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_2\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_1\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_3\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_2\ : std_logic;
signal \uart_tx.M_ctr_qZ1Z_4\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_3\ : std_logic;
signal \uart_tx.M_ctr_qZ1Z_5\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_5\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_4\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_5\ : std_logic;
signal \uart_tx.N_134_i\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \uart_tx.N_182_0\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_6\ : std_logic;
signal \uart_tx.N_143_0\ : std_logic;
signal \uart_tx.M_bitCtr_qZ0Z_1\ : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_4_cascade_\ : std_logic;
signal \uart_tx.M_bitCtr_qZ1Z_0\ : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_2\ : std_logic;
signal \uart_tx.M_txReg_d_3_7_ns_1_cascade_\ : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_1\ : std_logic;
signal \uart_tx.M_bitCtr_qZ0Z_2\ : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_5\ : std_logic;
signal btn_cond_out_16_5 : std_logic;
signal btn_cond_out_16_4 : std_logic;
signal btn_cond_out_17 : std_logic;
signal \click_dtct_M_last_q\ : std_logic;
signal \M_btn_cond_out_0_cascade_\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_0\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_1\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_2\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_3\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_4\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_5\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_6\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_7\ : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_8\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_9\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_10\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_11\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_12\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_13\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_14\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_15\ : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_16\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_17\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_18\ : std_logic;
signal \btn_cond.M_sync_out_i_g_0\ : std_logic;
signal \uart_tx.M_txReg_d_3\ : std_logic;
signal \uart_tx.M_state_qZ0Z_0\ : std_logic;
signal \uart_tx.M_state_qZ0Z_1\ : std_logic;
signal usb_tx_c : std_logic;
signal \uart_tx_N_186_1\ : std_logic;
signal \M_count_qZ0Z_0\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_0\ : std_logic;
signal \M_count_qZ0Z_6\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_6\ : std_logic;
signal \M_count_qZ0Z_4\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_4\ : std_logic;
signal \M_count_qZ0Z_7\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_7\ : std_logic;
signal \M_count_qZ0Z_2\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_2\ : std_logic;
signal \M_count_qZ0Z_3\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_3\ : std_logic;
signal \M_count_qZ0Z_1\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_1\ : std_logic;
signal \M_count_qZ0Z_5\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_5\ : std_logic;
signal \M_count_d6\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_6\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_5\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_4\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_7\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_11\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_8\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_10\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_9\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_15\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_14\ : std_logic;
signal \btn_cond.g0_13_cascade_\ : std_logic;
signal \btn_cond.g0_14\ : std_logic;
signal \btn_cond.g0_16_cascade_\ : std_logic;
signal \btn_cond.M_btn_cond_out_i_0\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_2\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_0\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_3\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_1\ : std_logic;
signal \btn_cond.g0_11\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_12\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_13\ : std_logic;
signal \btn_cond.g0_5\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_18\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_17\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_19\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_16\ : std_logic;
signal \btn_cond.g0_10\ : std_logic;
signal trigger_c : std_logic;
signal \btn_cond.sync.M_pipe_qZ0Z_0\ : std_logic;
signal clk_c_g : std_logic;
signal \btn_cond.sync.M_sync_out_0\ : std_logic;
signal \btn_cond.sync.M_sync_out_i_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal rst_n_wire : std_logic;
signal trigger_wire : std_logic;
signal usb_tx_wire : std_logic;

begin
    clk_wire <= clk;
    led <= led_wire;
    rst_n_wire <= rst_n;
    trigger_wire <= trigger;
    usb_tx <= usb_tx_wire;

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3296\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3298\,
            DIN => \N__3297\,
            DOUT => \N__3296\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3298\,
            PADOUT => \N__3297\,
            PADIN => \N__3296\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3287\,
            DIN => \N__3286\,
            DOUT => \N__3285\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3287\,
            PADOUT => \N__3286\,
            PADIN => \N__3285\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3278\,
            DIN => \N__3277\,
            DOUT => \N__3276\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3278\,
            PADOUT => \N__3277\,
            PADIN => \N__3276\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3269\,
            DIN => \N__3268\,
            DOUT => \N__3267\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3269\,
            PADOUT => \N__3268\,
            PADIN => \N__3267\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3260\,
            DIN => \N__3259\,
            DOUT => \N__3258\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3260\,
            PADOUT => \N__3259\,
            PADIN => \N__3258\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3251\,
            DIN => \N__3250\,
            DOUT => \N__3249\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3251\,
            PADOUT => \N__3250\,
            PADIN => \N__3249\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3242\,
            DIN => \N__3241\,
            DOUT => \N__3240\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3242\,
            PADOUT => \N__3241\,
            PADIN => \N__3240\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3233\,
            DIN => \N__3232\,
            DOUT => \N__3231\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3233\,
            PADOUT => \N__3232\,
            PADIN => \N__3231\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3224\,
            DIN => \N__3223\,
            DOUT => \N__3222\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3224\,
            PADOUT => \N__3223\,
            PADIN => \N__3222\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3215\,
            DIN => \N__3214\,
            DOUT => \N__3213\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3215\,
            PADOUT => \N__3214\,
            PADIN => \N__3213\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \trigger_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3206\,
            DIN => \N__3205\,
            DOUT => \N__3204\,
            PACKAGEPIN => trigger_wire
        );

    \trigger_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3206\,
            PADOUT => \N__3205\,
            PADIN => \N__3204\,
            CLOCKENABLE => 'H',
            DIN0 => trigger_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \usb_tx_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3197\,
            DIN => \N__3196\,
            DOUT => \N__3195\,
            PACKAGEPIN => usb_tx_wire
        );

    \usb_tx_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3197\,
            PADOUT => \N__3196\,
            PADIN => \N__3195\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2350\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__3178\,
            I => \btn_cond.g0_16_cascade_\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__3175\,
            I => \N__3171\
        );

    \I__713\ : InMux
    port map (
            O => \N__3174\,
            I => \N__3168\
        );

    \I__712\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3165\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3168\,
            I => \btn_cond.M_btn_cond_out_i_0\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3165\,
            I => \btn_cond.M_btn_cond_out_i_0\
        );

    \I__709\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3155\
        );

    \I__708\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3152\
        );

    \I__707\ : InMux
    port map (
            O => \N__3158\,
            I => \N__3149\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3155\,
            I => \N__3146\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3152\,
            I => \btn_cond.M_ctr_qZ0Z_2\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3149\,
            I => \btn_cond.M_ctr_qZ0Z_2\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__3146\,
            I => \btn_cond.M_ctr_qZ0Z_2\
        );

    \I__702\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3134\
        );

    \I__701\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3131\
        );

    \I__700\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3128\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3134\,
            I => \btn_cond.M_ctr_qZ0Z_0\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3131\,
            I => \btn_cond.M_ctr_qZ0Z_0\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3128\,
            I => \btn_cond.M_ctr_qZ0Z_0\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__3121\,
            I => \N__3116\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__3120\,
            I => \N__3113\
        );

    \I__694\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3110\
        );

    \I__693\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3107\
        );

    \I__692\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3104\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3110\,
            I => \btn_cond.M_ctr_qZ0Z_3\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3107\,
            I => \btn_cond.M_ctr_qZ0Z_3\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3104\,
            I => \btn_cond.M_ctr_qZ0Z_3\
        );

    \I__688\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3092\
        );

    \I__687\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3089\
        );

    \I__686\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3086\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3092\,
            I => \btn_cond.M_ctr_qZ0Z_1\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3089\,
            I => \btn_cond.M_ctr_qZ0Z_1\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3086\,
            I => \btn_cond.M_ctr_qZ0Z_1\
        );

    \I__682\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3076\,
            I => \btn_cond.g0_11\
        );

    \I__680\ : InMux
    port map (
            O => \N__3073\,
            I => \N__3068\
        );

    \I__679\ : InMux
    port map (
            O => \N__3072\,
            I => \N__3065\
        );

    \I__678\ : InMux
    port map (
            O => \N__3071\,
            I => \N__3062\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3068\,
            I => \btn_cond.M_ctr_qZ0Z_12\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3065\,
            I => \btn_cond.M_ctr_qZ0Z_12\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3062\,
            I => \btn_cond.M_ctr_qZ0Z_12\
        );

    \I__674\ : InMux
    port map (
            O => \N__3055\,
            I => \N__3052\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3052\,
            I => \N__3048\
        );

    \I__672\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3044\
        );

    \I__671\ : Span4Mux_v
    port map (
            O => \N__3048\,
            I => \N__3041\
        );

    \I__670\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3038\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3044\,
            I => \btn_cond.M_ctr_qZ0Z_13\
        );

    \I__668\ : Odrv4
    port map (
            O => \N__3041\,
            I => \btn_cond.M_ctr_qZ0Z_13\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3038\,
            I => \btn_cond.M_ctr_qZ0Z_13\
        );

    \I__666\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3028\,
            I => \btn_cond.g0_5\
        );

    \I__664\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3020\
        );

    \I__663\ : InMux
    port map (
            O => \N__3024\,
            I => \N__3017\
        );

    \I__662\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3014\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3020\,
            I => \btn_cond.M_ctr_qZ0Z_18\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3017\,
            I => \btn_cond.M_ctr_qZ0Z_18\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3014\,
            I => \btn_cond.M_ctr_qZ0Z_18\
        );

    \I__658\ : InMux
    port map (
            O => \N__3007\,
            I => \N__3003\
        );

    \I__657\ : InMux
    port map (
            O => \N__3006\,
            I => \N__2999\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3003\,
            I => \N__2996\
        );

    \I__655\ : InMux
    port map (
            O => \N__3002\,
            I => \N__2993\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__2999\,
            I => \btn_cond.M_ctr_qZ0Z_17\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__2996\,
            I => \btn_cond.M_ctr_qZ0Z_17\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__2993\,
            I => \btn_cond.M_ctr_qZ0Z_17\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__2986\,
            I => \N__2981\
        );

    \I__650\ : InMux
    port map (
            O => \N__2985\,
            I => \N__2978\
        );

    \I__649\ : InMux
    port map (
            O => \N__2984\,
            I => \N__2975\
        );

    \I__648\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2972\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__2978\,
            I => \btn_cond.M_ctr_qZ0Z_19\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__2975\,
            I => \btn_cond.M_ctr_qZ0Z_19\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__2972\,
            I => \btn_cond.M_ctr_qZ0Z_19\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__2965\,
            I => \N__2962\
        );

    \I__643\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2958\
        );

    \I__642\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2954\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__2958\,
            I => \N__2951\
        );

    \I__640\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2948\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__2954\,
            I => \btn_cond.M_ctr_qZ0Z_16\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__2951\,
            I => \btn_cond.M_ctr_qZ0Z_16\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__2948\,
            I => \btn_cond.M_ctr_qZ0Z_16\
        );

    \I__636\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2938\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__2938\,
            I => \btn_cond.g0_10\
        );

    \I__634\ : InMux
    port map (
            O => \N__2935\,
            I => \N__2932\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__2932\,
            I => \N__2929\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__2929\,
            I => \N__2926\
        );

    \I__631\ : Sp12to4
    port map (
            O => \N__2926\,
            I => \N__2923\
        );

    \I__630\ : Span12Mux_h
    port map (
            O => \N__2923\,
            I => \N__2920\
        );

    \I__629\ : Span12Mux_v
    port map (
            O => \N__2920\,
            I => \N__2917\
        );

    \I__628\ : Span12Mux_v
    port map (
            O => \N__2917\,
            I => \N__2914\
        );

    \I__627\ : Odrv12
    port map (
            O => \N__2914\,
            I => trigger_c
        );

    \I__626\ : InMux
    port map (
            O => \N__2911\,
            I => \N__2908\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__2908\,
            I => \btn_cond.sync.M_pipe_qZ0Z_0\
        );

    \I__624\ : ClkMux
    port map (
            O => \N__2905\,
            I => \N__2854\
        );

    \I__623\ : ClkMux
    port map (
            O => \N__2904\,
            I => \N__2854\
        );

    \I__622\ : ClkMux
    port map (
            O => \N__2903\,
            I => \N__2854\
        );

    \I__621\ : ClkMux
    port map (
            O => \N__2902\,
            I => \N__2854\
        );

    \I__620\ : ClkMux
    port map (
            O => \N__2901\,
            I => \N__2854\
        );

    \I__619\ : ClkMux
    port map (
            O => \N__2900\,
            I => \N__2854\
        );

    \I__618\ : ClkMux
    port map (
            O => \N__2899\,
            I => \N__2854\
        );

    \I__617\ : ClkMux
    port map (
            O => \N__2898\,
            I => \N__2854\
        );

    \I__616\ : ClkMux
    port map (
            O => \N__2897\,
            I => \N__2854\
        );

    \I__615\ : ClkMux
    port map (
            O => \N__2896\,
            I => \N__2854\
        );

    \I__614\ : ClkMux
    port map (
            O => \N__2895\,
            I => \N__2854\
        );

    \I__613\ : ClkMux
    port map (
            O => \N__2894\,
            I => \N__2854\
        );

    \I__612\ : ClkMux
    port map (
            O => \N__2893\,
            I => \N__2854\
        );

    \I__611\ : ClkMux
    port map (
            O => \N__2892\,
            I => \N__2854\
        );

    \I__610\ : ClkMux
    port map (
            O => \N__2891\,
            I => \N__2854\
        );

    \I__609\ : ClkMux
    port map (
            O => \N__2890\,
            I => \N__2854\
        );

    \I__608\ : ClkMux
    port map (
            O => \N__2889\,
            I => \N__2854\
        );

    \I__607\ : GlobalMux
    port map (
            O => \N__2854\,
            I => \N__2851\
        );

    \I__606\ : gio2CtrlBuf
    port map (
            O => \N__2851\,
            I => clk_c_g
        );

    \I__605\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__2845\,
            I => \btn_cond.sync.M_sync_out_0\
        );

    \I__603\ : IoInMux
    port map (
            O => \N__2842\,
            I => \N__2839\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__2839\,
            I => \btn_cond.sync.M_sync_out_i_0\
        );

    \I__601\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2833\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__2833\,
            I => \N__2830\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__2830\,
            I => \uart_tx.M_savedData_qZ0Z_7\
        );

    \I__598\ : InMux
    port map (
            O => \N__2827\,
            I => \N__2823\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__2826\,
            I => \N__2820\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__2823\,
            I => \N__2815\
        );

    \I__595\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2810\
        );

    \I__594\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2810\
        );

    \I__593\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2807\
        );

    \I__592\ : Odrv4
    port map (
            O => \N__2815\,
            I => \M_count_qZ0Z_2\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__2810\,
            I => \M_count_qZ0Z_2\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__2807\,
            I => \M_count_qZ0Z_2\
        );

    \I__589\ : InMux
    port map (
            O => \N__2800\,
            I => \N__2797\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__2797\,
            I => \uart_tx.M_savedData_qZ0Z_2\
        );

    \I__587\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2791\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__2791\,
            I => \N__2786\
        );

    \I__585\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2783\
        );

    \I__584\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2780\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__2786\,
            I => \M_count_qZ0Z_3\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__2783\,
            I => \M_count_qZ0Z_3\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__2780\,
            I => \M_count_qZ0Z_3\
        );

    \I__580\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2770\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__2770\,
            I => \uart_tx.M_savedData_qZ0Z_3\
        );

    \I__578\ : InMux
    port map (
            O => \N__2767\,
            I => \N__2762\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__2766\,
            I => \N__2759\
        );

    \I__576\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2756\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__2762\,
            I => \N__2752\
        );

    \I__574\ : InMux
    port map (
            O => \N__2759\,
            I => \N__2749\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__2756\,
            I => \N__2746\
        );

    \I__572\ : InMux
    port map (
            O => \N__2755\,
            I => \N__2743\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__2752\,
            I => \M_count_qZ0Z_1\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__2749\,
            I => \M_count_qZ0Z_1\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__2746\,
            I => \M_count_qZ0Z_1\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__2743\,
            I => \M_count_qZ0Z_1\
        );

    \I__567\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__2731\,
            I => \uart_tx.M_savedData_qZ0Z_1\
        );

    \I__565\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2725\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__2725\,
            I => \N__2720\
        );

    \I__563\ : InMux
    port map (
            O => \N__2724\,
            I => \N__2715\
        );

    \I__562\ : InMux
    port map (
            O => \N__2723\,
            I => \N__2715\
        );

    \I__561\ : Span4Mux_h
    port map (
            O => \N__2720\,
            I => \N__2709\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__2715\,
            I => \N__2709\
        );

    \I__559\ : InMux
    port map (
            O => \N__2714\,
            I => \N__2706\
        );

    \I__558\ : Odrv4
    port map (
            O => \N__2709\,
            I => \M_count_qZ0Z_5\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__2706\,
            I => \M_count_qZ0Z_5\
        );

    \I__556\ : InMux
    port map (
            O => \N__2701\,
            I => \N__2698\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__2698\,
            I => \uart_tx.M_savedData_qZ0Z_5\
        );

    \I__554\ : CEMux
    port map (
            O => \N__2695\,
            I => \N__2691\
        );

    \I__553\ : CEMux
    port map (
            O => \N__2694\,
            I => \N__2688\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__2691\,
            I => \M_count_d6\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__2688\,
            I => \M_count_d6\
        );

    \I__550\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2678\
        );

    \I__549\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2675\
        );

    \I__548\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2672\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__2678\,
            I => \btn_cond.M_ctr_qZ0Z_6\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2675\,
            I => \btn_cond.M_ctr_qZ0Z_6\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__2672\,
            I => \btn_cond.M_ctr_qZ0Z_6\
        );

    \I__544\ : InMux
    port map (
            O => \N__2665\,
            I => \N__2660\
        );

    \I__543\ : InMux
    port map (
            O => \N__2664\,
            I => \N__2657\
        );

    \I__542\ : InMux
    port map (
            O => \N__2663\,
            I => \N__2654\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__2660\,
            I => \btn_cond.M_ctr_qZ0Z_5\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2657\,
            I => \btn_cond.M_ctr_qZ0Z_5\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__2654\,
            I => \btn_cond.M_ctr_qZ0Z_5\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__2647\,
            I => \N__2642\
        );

    \I__537\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2639\
        );

    \I__536\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2636\
        );

    \I__535\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2633\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__2639\,
            I => \btn_cond.M_ctr_qZ0Z_4\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2636\,
            I => \btn_cond.M_ctr_qZ0Z_4\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2633\,
            I => \btn_cond.M_ctr_qZ0Z_4\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__2626\,
            I => \N__2623\
        );

    \I__530\ : InMux
    port map (
            O => \N__2623\,
            I => \N__2619\
        );

    \I__529\ : InMux
    port map (
            O => \N__2622\,
            I => \N__2615\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__2619\,
            I => \N__2612\
        );

    \I__527\ : InMux
    port map (
            O => \N__2618\,
            I => \N__2609\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__2615\,
            I => \btn_cond.M_ctr_qZ0Z_7\
        );

    \I__525\ : Odrv12
    port map (
            O => \N__2612\,
            I => \btn_cond.M_ctr_qZ0Z_7\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__2609\,
            I => \btn_cond.M_ctr_qZ0Z_7\
        );

    \I__523\ : InMux
    port map (
            O => \N__2602\,
            I => \N__2598\
        );

    \I__522\ : InMux
    port map (
            O => \N__2601\,
            I => \N__2594\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__2598\,
            I => \N__2591\
        );

    \I__520\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2588\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2594\,
            I => \btn_cond.M_ctr_qZ0Z_11\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__2591\,
            I => \btn_cond.M_ctr_qZ0Z_11\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__2588\,
            I => \btn_cond.M_ctr_qZ0Z_11\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__2581\,
            I => \N__2577\
        );

    \I__515\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2573\
        );

    \I__514\ : InMux
    port map (
            O => \N__2577\,
            I => \N__2570\
        );

    \I__513\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2567\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2573\,
            I => \btn_cond.M_ctr_qZ0Z_8\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__2570\,
            I => \btn_cond.M_ctr_qZ0Z_8\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__2567\,
            I => \btn_cond.M_ctr_qZ0Z_8\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__2560\,
            I => \N__2555\
        );

    \I__508\ : InMux
    port map (
            O => \N__2559\,
            I => \N__2552\
        );

    \I__507\ : InMux
    port map (
            O => \N__2558\,
            I => \N__2549\
        );

    \I__506\ : InMux
    port map (
            O => \N__2555\,
            I => \N__2546\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__2552\,
            I => \btn_cond.M_ctr_qZ0Z_10\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2549\,
            I => \btn_cond.M_ctr_qZ0Z_10\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2546\,
            I => \btn_cond.M_ctr_qZ0Z_10\
        );

    \I__502\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2534\
        );

    \I__501\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2531\
        );

    \I__500\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2528\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2534\,
            I => \btn_cond.M_ctr_qZ0Z_9\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__2531\,
            I => \btn_cond.M_ctr_qZ0Z_9\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2528\,
            I => \btn_cond.M_ctr_qZ0Z_9\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__2521\,
            I => \N__2517\
        );

    \I__495\ : InMux
    port map (
            O => \N__2520\,
            I => \N__2513\
        );

    \I__494\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2510\
        );

    \I__493\ : InMux
    port map (
            O => \N__2516\,
            I => \N__2507\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2513\,
            I => \btn_cond.M_ctr_qZ0Z_15\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2510\,
            I => \btn_cond.M_ctr_qZ0Z_15\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2507\,
            I => \btn_cond.M_ctr_qZ0Z_15\
        );

    \I__489\ : InMux
    port map (
            O => \N__2500\,
            I => \N__2495\
        );

    \I__488\ : InMux
    port map (
            O => \N__2499\,
            I => \N__2492\
        );

    \I__487\ : InMux
    port map (
            O => \N__2498\,
            I => \N__2489\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2495\,
            I => \btn_cond.M_ctr_qZ0Z_14\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__2492\,
            I => \btn_cond.M_ctr_qZ0Z_14\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__2489\,
            I => \btn_cond.M_ctr_qZ0Z_14\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__2482\,
            I => \btn_cond.g0_13_cascade_\
        );

    \I__482\ : InMux
    port map (
            O => \N__2479\,
            I => \N__2476\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2476\,
            I => \btn_cond.g0_14\
        );

    \I__480\ : InMux
    port map (
            O => \N__2473\,
            I => \bfn_15_27_0_\
        );

    \I__479\ : InMux
    port map (
            O => \N__2470\,
            I => \btn_cond.un1_M_ctr_q_cry_16\
        );

    \I__478\ : InMux
    port map (
            O => \N__2467\,
            I => \btn_cond.un1_M_ctr_q_cry_17\
        );

    \I__477\ : InMux
    port map (
            O => \N__2464\,
            I => \btn_cond.un1_M_ctr_q_cry_18\
        );

    \I__476\ : SRMux
    port map (
            O => \N__2461\,
            I => \N__2452\
        );

    \I__475\ : SRMux
    port map (
            O => \N__2460\,
            I => \N__2452\
        );

    \I__474\ : SRMux
    port map (
            O => \N__2459\,
            I => \N__2452\
        );

    \I__473\ : GlobalMux
    port map (
            O => \N__2452\,
            I => \N__2449\
        );

    \I__472\ : gio2CtrlBuf
    port map (
            O => \N__2449\,
            I => \btn_cond.M_sync_out_i_g_0\
        );

    \I__471\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2443\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2443\,
            I => \uart_tx.M_txReg_d_3\
        );

    \I__469\ : InMux
    port map (
            O => \N__2440\,
            I => \N__2437\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2437\,
            I => \N__2430\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__2436\,
            I => \N__2427\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__2435\,
            I => \N__2421\
        );

    \I__465\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2415\
        );

    \I__464\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2415\
        );

    \I__463\ : Span4Mux_h
    port map (
            O => \N__2430\,
            I => \N__2412\
        );

    \I__462\ : InMux
    port map (
            O => \N__2427\,
            I => \N__2403\
        );

    \I__461\ : InMux
    port map (
            O => \N__2426\,
            I => \N__2403\
        );

    \I__460\ : InMux
    port map (
            O => \N__2425\,
            I => \N__2403\
        );

    \I__459\ : InMux
    port map (
            O => \N__2424\,
            I => \N__2403\
        );

    \I__458\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2398\
        );

    \I__457\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2398\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2415\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__2412\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2403\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2398\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__452\ : InMux
    port map (
            O => \N__2389\,
            I => \N__2385\
        );

    \I__451\ : CascadeMux
    port map (
            O => \N__2388\,
            I => \N__2379\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2385\,
            I => \N__2373\
        );

    \I__449\ : InMux
    port map (
            O => \N__2384\,
            I => \N__2366\
        );

    \I__448\ : InMux
    port map (
            O => \N__2383\,
            I => \N__2366\
        );

    \I__447\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2366\
        );

    \I__446\ : InMux
    port map (
            O => \N__2379\,
            I => \N__2357\
        );

    \I__445\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2357\
        );

    \I__444\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2357\
        );

    \I__443\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2357\
        );

    \I__442\ : Odrv4
    port map (
            O => \N__2373\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2366\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2357\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__439\ : IoInMux
    port map (
            O => \N__2350\,
            I => \N__2347\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2347\,
            I => \N__2344\
        );

    \I__437\ : Span4Mux_s0_v
    port map (
            O => \N__2344\,
            I => \N__2341\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__2341\,
            I => \N__2338\
        );

    \I__435\ : Span12Mux_h
    port map (
            O => \N__2338\,
            I => \N__2335\
        );

    \I__434\ : Span12Mux_v
    port map (
            O => \N__2335\,
            I => \N__2332\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__2332\,
            I => usb_tx_c
        );

    \I__432\ : SRMux
    port map (
            O => \N__2329\,
            I => \N__2324\
        );

    \I__431\ : InMux
    port map (
            O => \N__2328\,
            I => \N__2318\
        );

    \I__430\ : InMux
    port map (
            O => \N__2327\,
            I => \N__2318\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2324\,
            I => \N__2306\
        );

    \I__428\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2300\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2318\,
            I => \N__2297\
        );

    \I__426\ : InMux
    port map (
            O => \N__2317\,
            I => \N__2294\
        );

    \I__425\ : InMux
    port map (
            O => \N__2316\,
            I => \N__2287\
        );

    \I__424\ : InMux
    port map (
            O => \N__2315\,
            I => \N__2287\
        );

    \I__423\ : InMux
    port map (
            O => \N__2314\,
            I => \N__2287\
        );

    \I__422\ : InMux
    port map (
            O => \N__2313\,
            I => \N__2282\
        );

    \I__421\ : InMux
    port map (
            O => \N__2312\,
            I => \N__2282\
        );

    \I__420\ : InMux
    port map (
            O => \N__2311\,
            I => \N__2275\
        );

    \I__419\ : InMux
    port map (
            O => \N__2310\,
            I => \N__2275\
        );

    \I__418\ : InMux
    port map (
            O => \N__2309\,
            I => \N__2275\
        );

    \I__417\ : Span4Mux_h
    port map (
            O => \N__2306\,
            I => \N__2272\
        );

    \I__416\ : InMux
    port map (
            O => \N__2305\,
            I => \N__2269\
        );

    \I__415\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2266\
        );

    \I__414\ : InMux
    port map (
            O => \N__2303\,
            I => \N__2263\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2300\,
            I => \uart_tx_N_186_1\
        );

    \I__412\ : Odrv4
    port map (
            O => \N__2297\,
            I => \uart_tx_N_186_1\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2294\,
            I => \uart_tx_N_186_1\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2287\,
            I => \uart_tx_N_186_1\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2282\,
            I => \uart_tx_N_186_1\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2275\,
            I => \uart_tx_N_186_1\
        );

    \I__407\ : Odrv4
    port map (
            O => \N__2272\,
            I => \uart_tx_N_186_1\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2269\,
            I => \uart_tx_N_186_1\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2266\,
            I => \uart_tx_N_186_1\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2263\,
            I => \uart_tx_N_186_1\
        );

    \I__403\ : InMux
    port map (
            O => \N__2242\,
            I => \N__2239\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2239\,
            I => \N__2235\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__2238\,
            I => \N__2231\
        );

    \I__400\ : Span4Mux_v
    port map (
            O => \N__2235\,
            I => \N__2227\
        );

    \I__399\ : InMux
    port map (
            O => \N__2234\,
            I => \N__2224\
        );

    \I__398\ : InMux
    port map (
            O => \N__2231\,
            I => \N__2219\
        );

    \I__397\ : InMux
    port map (
            O => \N__2230\,
            I => \N__2219\
        );

    \I__396\ : Odrv4
    port map (
            O => \N__2227\,
            I => \M_count_qZ0Z_0\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2224\,
            I => \M_count_qZ0Z_0\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2219\,
            I => \M_count_qZ0Z_0\
        );

    \I__393\ : InMux
    port map (
            O => \N__2212\,
            I => \N__2209\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2209\,
            I => \N__2206\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__2206\,
            I => \uart_tx.M_savedData_qZ0Z_0\
        );

    \I__390\ : InMux
    port map (
            O => \N__2203\,
            I => \N__2200\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2200\,
            I => \N__2195\
        );

    \I__388\ : InMux
    port map (
            O => \N__2199\,
            I => \N__2192\
        );

    \I__387\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2189\
        );

    \I__386\ : Span4Mux_v
    port map (
            O => \N__2195\,
            I => \N__2184\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2192\,
            I => \N__2184\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2189\,
            I => \N__2181\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__2184\,
            I => \M_count_qZ0Z_6\
        );

    \I__382\ : Odrv4
    port map (
            O => \N__2181\,
            I => \M_count_qZ0Z_6\
        );

    \I__381\ : InMux
    port map (
            O => \N__2176\,
            I => \N__2173\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2173\,
            I => \uart_tx.M_savedData_qZ0Z_6\
        );

    \I__379\ : InMux
    port map (
            O => \N__2170\,
            I => \N__2167\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2167\,
            I => \N__2164\
        );

    \I__377\ : Span4Mux_h
    port map (
            O => \N__2164\,
            I => \N__2159\
        );

    \I__376\ : InMux
    port map (
            O => \N__2163\,
            I => \N__2156\
        );

    \I__375\ : InMux
    port map (
            O => \N__2162\,
            I => \N__2153\
        );

    \I__374\ : Odrv4
    port map (
            O => \N__2159\,
            I => \M_count_qZ0Z_4\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2156\,
            I => \M_count_qZ0Z_4\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2153\,
            I => \M_count_qZ0Z_4\
        );

    \I__371\ : InMux
    port map (
            O => \N__2146\,
            I => \N__2143\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2143\,
            I => \uart_tx.M_savedData_qZ0Z_4\
        );

    \I__369\ : InMux
    port map (
            O => \N__2140\,
            I => \N__2137\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2137\,
            I => \N__2134\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__2134\,
            I => \N__2130\
        );

    \I__366\ : InMux
    port map (
            O => \N__2133\,
            I => \N__2127\
        );

    \I__365\ : Odrv4
    port map (
            O => \N__2130\,
            I => \M_count_qZ0Z_7\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2127\,
            I => \M_count_qZ0Z_7\
        );

    \I__363\ : InMux
    port map (
            O => \N__2122\,
            I => \btn_cond.un1_M_ctr_q_cry_6\
        );

    \I__362\ : InMux
    port map (
            O => \N__2119\,
            I => \bfn_15_26_0_\
        );

    \I__361\ : InMux
    port map (
            O => \N__2116\,
            I => \btn_cond.un1_M_ctr_q_cry_8\
        );

    \I__360\ : InMux
    port map (
            O => \N__2113\,
            I => \btn_cond.un1_M_ctr_q_cry_9\
        );

    \I__359\ : InMux
    port map (
            O => \N__2110\,
            I => \btn_cond.un1_M_ctr_q_cry_10\
        );

    \I__358\ : InMux
    port map (
            O => \N__2107\,
            I => \btn_cond.un1_M_ctr_q_cry_11\
        );

    \I__357\ : InMux
    port map (
            O => \N__2104\,
            I => \btn_cond.un1_M_ctr_q_cry_12\
        );

    \I__356\ : InMux
    port map (
            O => \N__2101\,
            I => \btn_cond.un1_M_ctr_q_cry_13\
        );

    \I__355\ : InMux
    port map (
            O => \N__2098\,
            I => \btn_cond.un1_M_ctr_q_cry_14\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2095\,
            I => \N__2092\
        );

    \I__353\ : InMux
    port map (
            O => \N__2092\,
            I => \N__2083\
        );

    \I__352\ : InMux
    port map (
            O => \N__2091\,
            I => \N__2083\
        );

    \I__351\ : InMux
    port map (
            O => \N__2090\,
            I => \N__2080\
        );

    \I__350\ : InMux
    port map (
            O => \N__2089\,
            I => \N__2077\
        );

    \I__349\ : InMux
    port map (
            O => \N__2088\,
            I => \N__2074\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2083\,
            I => btn_cond_out_16_5
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2080\,
            I => btn_cond_out_16_5
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2077\,
            I => btn_cond_out_16_5
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2074\,
            I => btn_cond_out_16_5
        );

    \I__344\ : InMux
    port map (
            O => \N__2065\,
            I => \N__2058\
        );

    \I__343\ : InMux
    port map (
            O => \N__2064\,
            I => \N__2055\
        );

    \I__342\ : InMux
    port map (
            O => \N__2063\,
            I => \N__2050\
        );

    \I__341\ : InMux
    port map (
            O => \N__2062\,
            I => \N__2050\
        );

    \I__340\ : InMux
    port map (
            O => \N__2061\,
            I => \N__2047\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2058\,
            I => \N__2044\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2055\,
            I => \N__2041\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2050\,
            I => btn_cond_out_16_4
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2047\,
            I => btn_cond_out_16_4
        );

    \I__335\ : Odrv4
    port map (
            O => \N__2044\,
            I => btn_cond_out_16_4
        );

    \I__334\ : Odrv4
    port map (
            O => \N__2041\,
            I => btn_cond_out_16_4
        );

    \I__333\ : InMux
    port map (
            O => \N__2032\,
            I => \N__2026\
        );

    \I__332\ : InMux
    port map (
            O => \N__2031\,
            I => \N__2023\
        );

    \I__331\ : InMux
    port map (
            O => \N__2030\,
            I => \N__2020\
        );

    \I__330\ : InMux
    port map (
            O => \N__2029\,
            I => \N__2017\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2026\,
            I => btn_cond_out_17
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2023\,
            I => btn_cond_out_17
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2020\,
            I => btn_cond_out_17
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2017\,
            I => btn_cond_out_17
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2008\,
            I => \N__2001\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2007\,
            I => \N__1998\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__2006\,
            I => \N__1994\
        );

    \I__322\ : InMux
    port map (
            O => \N__2005\,
            I => \N__1991\
        );

    \I__321\ : InMux
    port map (
            O => \N__2004\,
            I => \N__1988\
        );

    \I__320\ : InMux
    port map (
            O => \N__2001\,
            I => \N__1985\
        );

    \I__319\ : InMux
    port map (
            O => \N__1998\,
            I => \N__1982\
        );

    \I__318\ : InMux
    port map (
            O => \N__1997\,
            I => \N__1977\
        );

    \I__317\ : InMux
    port map (
            O => \N__1994\,
            I => \N__1977\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1991\,
            I => \click_dtct_M_last_q\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__1988\,
            I => \click_dtct_M_last_q\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__1985\,
            I => \click_dtct_M_last_q\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__1982\,
            I => \click_dtct_M_last_q\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__1977\,
            I => \click_dtct_M_last_q\
        );

    \I__311\ : CascadeMux
    port map (
            O => \N__1966\,
            I => \M_btn_cond_out_0_cascade_\
        );

    \I__310\ : InMux
    port map (
            O => \N__1963\,
            I => \btn_cond.un1_M_ctr_q_cry_0\
        );

    \I__309\ : InMux
    port map (
            O => \N__1960\,
            I => \btn_cond.un1_M_ctr_q_cry_1\
        );

    \I__308\ : InMux
    port map (
            O => \N__1957\,
            I => \btn_cond.un1_M_ctr_q_cry_2\
        );

    \I__307\ : InMux
    port map (
            O => \N__1954\,
            I => \btn_cond.un1_M_ctr_q_cry_3\
        );

    \I__306\ : InMux
    port map (
            O => \N__1951\,
            I => \btn_cond.un1_M_ctr_q_cry_4\
        );

    \I__305\ : InMux
    port map (
            O => \N__1948\,
            I => \btn_cond.un1_M_ctr_q_cry_5\
        );

    \I__304\ : InMux
    port map (
            O => \N__1945\,
            I => \uart_tx.un1_M_ctr_q_3_cry_5\
        );

    \I__303\ : CascadeMux
    port map (
            O => \N__1942\,
            I => \N__1938\
        );

    \I__302\ : InMux
    port map (
            O => \N__1941\,
            I => \N__1935\
        );

    \I__301\ : InMux
    port map (
            O => \N__1938\,
            I => \N__1932\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1935\,
            I => \uart_tx.N_134_i\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1932\,
            I => \uart_tx.N_134_i\
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__1927\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\
        );

    \I__297\ : InMux
    port map (
            O => \N__1924\,
            I => \N__1915\
        );

    \I__296\ : InMux
    port map (
            O => \N__1923\,
            I => \N__1908\
        );

    \I__295\ : InMux
    port map (
            O => \N__1922\,
            I => \N__1908\
        );

    \I__294\ : InMux
    port map (
            O => \N__1921\,
            I => \N__1908\
        );

    \I__293\ : InMux
    port map (
            O => \N__1920\,
            I => \N__1901\
        );

    \I__292\ : InMux
    port map (
            O => \N__1919\,
            I => \N__1901\
        );

    \I__291\ : InMux
    port map (
            O => \N__1918\,
            I => \N__1901\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1915\,
            I => \uart_tx.N_182_0\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__1908\,
            I => \uart_tx.N_182_0\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1901\,
            I => \uart_tx.N_182_0\
        );

    \I__287\ : InMux
    port map (
            O => \N__1894\,
            I => \N__1890\
        );

    \I__286\ : InMux
    port map (
            O => \N__1893\,
            I => \N__1887\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__1890\,
            I => \uart_tx.M_ctr_qZ0Z_6\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1887\,
            I => \uart_tx.M_ctr_qZ0Z_6\
        );

    \I__283\ : CascadeMux
    port map (
            O => \N__1882\,
            I => \N__1879\
        );

    \I__282\ : InMux
    port map (
            O => \N__1879\,
            I => \N__1876\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__1876\,
            I => \uart_tx.N_143_0\
        );

    \I__280\ : InMux
    port map (
            O => \N__1873\,
            I => \N__1865\
        );

    \I__279\ : InMux
    port map (
            O => \N__1872\,
            I => \N__1865\
        );

    \I__278\ : InMux
    port map (
            O => \N__1871\,
            I => \N__1860\
        );

    \I__277\ : InMux
    port map (
            O => \N__1870\,
            I => \N__1860\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1865\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1860\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__1855\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_4_cascade_\
        );

    \I__273\ : InMux
    port map (
            O => \N__1852\,
            I => \N__1849\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1849\,
            I => \N__1842\
        );

    \I__271\ : InMux
    port map (
            O => \N__1848\,
            I => \N__1839\
        );

    \I__270\ : InMux
    port map (
            O => \N__1847\,
            I => \N__1834\
        );

    \I__269\ : InMux
    port map (
            O => \N__1846\,
            I => \N__1834\
        );

    \I__268\ : InMux
    port map (
            O => \N__1845\,
            I => \N__1831\
        );

    \I__267\ : Odrv4
    port map (
            O => \N__1842\,
            I => \uart_tx.M_bitCtr_qZ1Z_0\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1839\,
            I => \uart_tx.M_bitCtr_qZ1Z_0\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1834\,
            I => \uart_tx.M_bitCtr_qZ1Z_0\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1831\,
            I => \uart_tx.M_bitCtr_qZ1Z_0\
        );

    \I__263\ : InMux
    port map (
            O => \N__1822\,
            I => \N__1819\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1819\,
            I => \N__1816\
        );

    \I__261\ : Odrv4
    port map (
            O => \N__1816\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_2\
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__1813\,
            I => \uart_tx.M_txReg_d_3_7_ns_1_cascade_\
        );

    \I__259\ : InMux
    port map (
            O => \N__1810\,
            I => \N__1807\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__1807\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_1\
        );

    \I__257\ : InMux
    port map (
            O => \N__1804\,
            I => \N__1796\
        );

    \I__256\ : InMux
    port map (
            O => \N__1803\,
            I => \N__1785\
        );

    \I__255\ : InMux
    port map (
            O => \N__1802\,
            I => \N__1785\
        );

    \I__254\ : InMux
    port map (
            O => \N__1801\,
            I => \N__1785\
        );

    \I__253\ : InMux
    port map (
            O => \N__1800\,
            I => \N__1785\
        );

    \I__252\ : InMux
    port map (
            O => \N__1799\,
            I => \N__1785\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1796\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1785\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__249\ : InMux
    port map (
            O => \N__1780\,
            I => \N__1777\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1777\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_5\
        );

    \I__247\ : InMux
    port map (
            O => \N__1774\,
            I => \N__1771\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1771\,
            I => \reset_cond.M_stage_qZ0Z_2\
        );

    \I__245\ : InMux
    port map (
            O => \N__1768\,
            I => \N__1765\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1765\,
            I => \N__1759\
        );

    \I__243\ : InMux
    port map (
            O => \N__1764\,
            I => \N__1752\
        );

    \I__242\ : InMux
    port map (
            O => \N__1763\,
            I => \N__1752\
        );

    \I__241\ : InMux
    port map (
            O => \N__1762\,
            I => \N__1752\
        );

    \I__240\ : Span4Mux_h
    port map (
            O => \N__1759\,
            I => \N__1749\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1752\,
            I => \N__1746\
        );

    \I__238\ : Sp12to4
    port map (
            O => \N__1749\,
            I => \N__1741\
        );

    \I__237\ : Span12Mux_h
    port map (
            O => \N__1746\,
            I => \N__1741\
        );

    \I__236\ : Span12Mux_v
    port map (
            O => \N__1741\,
            I => \N__1738\
        );

    \I__235\ : Odrv12
    port map (
            O => \N__1738\,
            I => rst_n_c
        );

    \I__234\ : InMux
    port map (
            O => \N__1735\,
            I => \N__1732\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1732\,
            I => \reset_cond.M_stage_qZ0Z_0\
        );

    \I__232\ : InMux
    port map (
            O => \N__1729\,
            I => \N__1726\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1726\,
            I => \reset_cond.M_stage_qZ0Z_1\
        );

    \I__230\ : CascadeMux
    port map (
            O => \N__1723\,
            I => \N__1719\
        );

    \I__229\ : InMux
    port map (
            O => \N__1722\,
            I => \N__1716\
        );

    \I__228\ : InMux
    port map (
            O => \N__1719\,
            I => \N__1713\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__1716\,
            I => \uart_tx.N_186_1_i\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1713\,
            I => \uart_tx.N_186_1_i\
        );

    \I__225\ : InMux
    port map (
            O => \N__1708\,
            I => \N__1704\
        );

    \I__224\ : InMux
    port map (
            O => \N__1707\,
            I => \N__1701\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1704\,
            I => \uart_tx.M_ctr_qZ0Z_0\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1701\,
            I => \uart_tx.M_ctr_qZ0Z_0\
        );

    \I__221\ : CascadeMux
    port map (
            O => \N__1696\,
            I => \N__1692\
        );

    \I__220\ : InMux
    port map (
            O => \N__1695\,
            I => \N__1689\
        );

    \I__219\ : InMux
    port map (
            O => \N__1692\,
            I => \N__1686\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1689\,
            I => \uart_tx.M_ctr_qZ1Z_1\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1686\,
            I => \uart_tx.M_ctr_qZ1Z_1\
        );

    \I__216\ : InMux
    port map (
            O => \N__1681\,
            I => \uart_tx.un1_M_ctr_q_3_cry_0\
        );

    \I__215\ : InMux
    port map (
            O => \N__1678\,
            I => \N__1674\
        );

    \I__214\ : InMux
    port map (
            O => \N__1677\,
            I => \N__1671\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1674\,
            I => \uart_tx.M_ctr_qZ0Z_2\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1671\,
            I => \uart_tx.M_ctr_qZ0Z_2\
        );

    \I__211\ : InMux
    port map (
            O => \N__1666\,
            I => \N__1663\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1663\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_2\
        );

    \I__209\ : InMux
    port map (
            O => \N__1660\,
            I => \uart_tx.un1_M_ctr_q_3_cry_1\
        );

    \I__208\ : InMux
    port map (
            O => \N__1657\,
            I => \N__1653\
        );

    \I__207\ : InMux
    port map (
            O => \N__1656\,
            I => \N__1650\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1653\,
            I => \uart_tx.M_ctr_qZ0Z_3\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__1650\,
            I => \uart_tx.M_ctr_qZ0Z_3\
        );

    \I__204\ : InMux
    port map (
            O => \N__1645\,
            I => \uart_tx.un1_M_ctr_q_3_cry_2\
        );

    \I__203\ : InMux
    port map (
            O => \N__1642\,
            I => \N__1638\
        );

    \I__202\ : InMux
    port map (
            O => \N__1641\,
            I => \N__1635\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1638\,
            I => \uart_tx.M_ctr_qZ1Z_4\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1635\,
            I => \uart_tx.M_ctr_qZ1Z_4\
        );

    \I__199\ : InMux
    port map (
            O => \N__1630\,
            I => \uart_tx.un1_M_ctr_q_3_cry_3\
        );

    \I__198\ : InMux
    port map (
            O => \N__1627\,
            I => \N__1623\
        );

    \I__197\ : InMux
    port map (
            O => \N__1626\,
            I => \N__1620\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1623\,
            I => \uart_tx.M_ctr_qZ1Z_5\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1620\,
            I => \uart_tx.M_ctr_qZ1Z_5\
        );

    \I__194\ : InMux
    port map (
            O => \N__1615\,
            I => \N__1612\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1612\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_5\
        );

    \I__192\ : InMux
    port map (
            O => \N__1609\,
            I => \uart_tx.un1_M_ctr_q_3_cry_4\
        );

    \I__191\ : InMux
    port map (
            O => \N__1606\,
            I => \N__1603\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1603\,
            I => \un1_M_count_q_axbxc7_1\
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__1600\,
            I => \btn_cond.out_17_6_cascade_\
        );

    \I__188\ : InMux
    port map (
            O => \N__1597\,
            I => \N__1594\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1594\,
            I => \btn_cond.out_17_8\
        );

    \I__186\ : CascadeMux
    port map (
            O => \N__1591\,
            I => \btn_cond_out_17_cascade_\
        );

    \I__185\ : InMux
    port map (
            O => \N__1588\,
            I => \N__1582\
        );

    \I__184\ : InMux
    port map (
            O => \N__1587\,
            I => \N__1575\
        );

    \I__183\ : InMux
    port map (
            O => \N__1586\,
            I => \N__1575\
        );

    \I__182\ : InMux
    port map (
            O => \N__1585\,
            I => \N__1575\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1582\,
            I => \N__1572\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1575\,
            I => click_dtct_out8
        );

    \I__179\ : Odrv4
    port map (
            O => \N__1572\,
            I => click_dtct_out8
        );

    \I__178\ : InMux
    port map (
            O => \N__1567\,
            I => \N__1564\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1564\,
            I => \btn_cond.out_17_7\
        );

    \I__176\ : CascadeMux
    port map (
            O => \N__1561\,
            I => \click_dtct_M_count_d6_0_1_cascade_\
        );

    \I__175\ : CascadeMux
    port map (
            O => \N__1558\,
            I => \uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_\
        );

    \I__174\ : InMux
    port map (
            O => \N__1555\,
            I => \N__1552\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1552\,
            I => \uart_tx_N_187\
        );

    \I__172\ : CascadeMux
    port map (
            O => \N__1549\,
            I => \un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_\
        );

    \I__171\ : InMux
    port map (
            O => \N__1546\,
            I => \N__1543\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1543\,
            I => \un1_M_count_q_ac0_5_m2_0_a2_3\
        );

    \I__169\ : CascadeMux
    port map (
            O => \N__1540\,
            I => \un1_M_count_q_ac0_5_m2_0_a2_3_cascade_\
        );

    \I__168\ : InMux
    port map (
            O => \N__1537\,
            I => \N__1533\
        );

    \I__167\ : InMux
    port map (
            O => \N__1536\,
            I => \N__1530\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1533\,
            I => \un1_M_count_q_ac0_out\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1530\,
            I => \un1_M_count_q_ac0_out\
        );

    \I__164\ : InMux
    port map (
            O => \N__1525\,
            I => \N__1516\
        );

    \I__163\ : InMux
    port map (
            O => \N__1524\,
            I => \N__1516\
        );

    \I__162\ : InMux
    port map (
            O => \N__1523\,
            I => \N__1513\
        );

    \I__161\ : InMux
    port map (
            O => \N__1522\,
            I => \N__1510\
        );

    \I__160\ : InMux
    port map (
            O => \N__1521\,
            I => \N__1507\
        );

    \I__159\ : LocalMux
    port map (
            O => \N__1516\,
            I => click_dtct_out3
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1513\,
            I => click_dtct_out3
        );

    \I__157\ : LocalMux
    port map (
            O => \N__1510\,
            I => click_dtct_out3
        );

    \I__156\ : LocalMux
    port map (
            O => \N__1507\,
            I => click_dtct_out3
        );

    \I__155\ : SRMux
    port map (
            O => \N__1498\,
            I => \N__1493\
        );

    \I__154\ : SRMux
    port map (
            O => \N__1497\,
            I => \N__1490\
        );

    \I__153\ : SRMux
    port map (
            O => \N__1496\,
            I => \N__1487\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1493\,
            I => \N__1484\
        );

    \I__151\ : LocalMux
    port map (
            O => \N__1490\,
            I => \N__1480\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1487\,
            I => \N__1477\
        );

    \I__149\ : Span4Mux_v
    port map (
            O => \N__1484\,
            I => \N__1474\
        );

    \I__148\ : InMux
    port map (
            O => \N__1483\,
            I => \N__1471\
        );

    \I__147\ : Span4Mux_v
    port map (
            O => \N__1480\,
            I => \N__1467\
        );

    \I__146\ : Span4Mux_v
    port map (
            O => \N__1477\,
            I => \N__1460\
        );

    \I__145\ : Span4Mux_h
    port map (
            O => \N__1474\,
            I => \N__1460\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__1471\,
            I => \N__1460\
        );

    \I__143\ : InMux
    port map (
            O => \N__1470\,
            I => \N__1457\
        );

    \I__142\ : Odrv4
    port map (
            O => \N__1467\,
            I => \M_reset_cond_out_0\
        );

    \I__141\ : Odrv4
    port map (
            O => \N__1460\,
            I => \M_reset_cond_out_0\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1457\,
            I => \M_reset_cond_out_0\
        );

    \I__139\ : CascadeMux
    port map (
            O => \N__1450\,
            I => \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\
        );

    \I__138\ : CascadeMux
    port map (
            O => \N__1447\,
            I => \uart_tx.N_182_0_cascade_\
        );

    \I__137\ : CascadeMux
    port map (
            O => \N__1444\,
            I => \uart_tx.N_143_0_cascade_\
        );

    \I__136\ : CascadeMux
    port map (
            O => \N__1441\,
            I => \uart_tx_N_185_cascade_\
        );

    \I__135\ : InMux
    port map (
            O => \N__1438\,
            I => \N__1435\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__1435\,
            I => \un1_M_count_q_ac0_1\
        );

    \I__133\ : CascadeMux
    port map (
            O => \N__1432\,
            I => \click_dtct_out3_cascade_\
        );

    \I__132\ : CascadeMux
    port map (
            O => \N__1429\,
            I => \un1_M_count_q_ac0_7_cascade_\
        );

    \I__131\ : InMux
    port map (
            O => \N__1426\,
            I => \N__1414\
        );

    \I__130\ : InMux
    port map (
            O => \N__1425\,
            I => \N__1414\
        );

    \I__129\ : InMux
    port map (
            O => \N__1424\,
            I => \N__1414\
        );

    \I__128\ : InMux
    port map (
            O => \N__1423\,
            I => \N__1414\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1414\,
            I => click_dtct_out_d
        );

    \I__126\ : CascadeMux
    port map (
            O => \N__1411\,
            I => \click_dtct_out_d_cascade_\
        );

    \I__125\ : InMux
    port map (
            O => \N__1408\,
            I => \N__1404\
        );

    \I__124\ : InMux
    port map (
            O => \N__1407\,
            I => \N__1401\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1404\,
            I => \un1_M_count_q_ac0_7\
        );

    \I__122\ : LocalMux
    port map (
            O => \N__1401\,
            I => \un1_M_count_q_ac0_7\
        );

    \I__121\ : CascadeMux
    port map (
            O => \N__1396\,
            I => \uart_tx.N_134_i_cascade_\
        );

    \I__120\ : CascadeMux
    port map (
            O => \N__1393\,
            I => \un1_M_count_q_ac0_1_cascade_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \btn_cond.un1_M_ctr_q_cry_7\,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \btn_cond.un1_M_ctr_q_cry_15\,
            carryinitout => \bfn_15_27_0_\
        );

    \btn_cond.sync.M_pipe_q_RNIJLM5_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2842\,
            GLOBALBUFFEROUTPUT => \btn_cond.M_sync_out_i_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \M_count_q_RNI2B741_0_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2234\,
            in2 => \_gnd_net_\,
            in3 => \N__2303\,
            lcout => \un1_M_count_q_ac0_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNI0H5P2_1_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__2765\,
            in1 => \N__1536\,
            in2 => \N__2008\,
            in3 => \N__1521\,
            lcout => \un1_M_count_q_ac0_1\,
            ltout => \un1_M_count_q_ac0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_2_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2819\,
            in2 => \N__1393\,
            in3 => \N__1423\,
            lcout => \M_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2900\,
            ce => 'H',
            sr => \N__1498\
        );

    \M_count_q_5_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__2723\,
            in1 => \N__1424\,
            in2 => \_gnd_net_\,
            in3 => \N__1407\,
            lcout => \M_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2900\,
            ce => 'H',
            sr => \N__1498\
        );

    \M_count_q_3_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__1425\,
            in1 => \N__2790\,
            in2 => \N__2826\,
            in3 => \N__1438\,
            lcout => \M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2900\,
            ce => 'H',
            sr => \N__1498\
        );

    \click_dtct.M_last_q_RNIUTK51_1_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2088\,
            in1 => \N__2064\,
            in2 => \N__2006\,
            in3 => \N__2029\,
            lcout => click_dtct_out3,
            ltout => \click_dtct_out3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIGFD24_4_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__1546\,
            in1 => \N__2162\,
            in2 => \N__1432\,
            in3 => \N__1997\,
            lcout => \un1_M_count_q_ac0_7\,
            ltout => \un1_M_count_q_ac0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_6_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__2724\,
            in1 => \N__2199\,
            in2 => \N__1429\,
            in3 => \N__1426\,
            lcout => \M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2900\,
            ce => 'H',
            sr => \N__1498\
        );

    \click_dtct.M_last_q_RNIUTK51_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__2090\,
            in1 => \N__2061\,
            in2 => \N__2007\,
            in3 => \N__2031\,
            lcout => click_dtct_out_d,
            ltout => \click_dtct_out_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_7_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101010101010"
        )
    port map (
            in0 => \N__2133\,
            in1 => \N__1606\,
            in2 => \N__1411\,
            in3 => \N__1408\,
            lcout => \M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2903\,
            ce => 'H',
            sr => \N__1496\
        );

    \reset_cond.M_stage_q_3_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1768\,
            in2 => \_gnd_net_\,
            in3 => \N__1774\,
            lcout => \M_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2892\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_5_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__2313\,
            in1 => \N__1615\,
            in2 => \N__1942\,
            in3 => \N__1922\,
            lcout => \uart_tx.M_ctr_qZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_0_1_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__2377\,
            in1 => \_gnd_net_\,
            in2 => \N__2435\,
            in3 => \_gnd_net_\,
            lcout => \uart_tx.N_134_i\,
            ltout => \uart_tx.N_134_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_2_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__2312\,
            in1 => \N__1666\,
            in2 => \N__1396\,
            in3 => \N__1921\,
            lcout => \uart_tx.M_ctr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_1_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__1923\,
            in1 => \N__1470\,
            in2 => \N__2388\,
            in3 => \N__2434\,
            lcout => \uart_tx.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_1_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2420\,
            in2 => \_gnd_net_\,
            in3 => \N__2376\,
            lcout => \uart_tx.N_186_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNIGGUF1_0_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__1626\,
            in1 => \N__1677\,
            in2 => \N__1696\,
            in3 => \N__1707\,
            lcout => OPEN,
            ltout => \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNI3KTJ2_6_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__1893\,
            in1 => \N__1641\,
            in2 => \N__1450\,
            in3 => \N__1656\,
            lcout => \uart_tx.N_182_0\,
            ltout => \uart_tx.N_182_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_0_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000101000"
        )
    port map (
            in0 => \N__2378\,
            in1 => \N__1852\,
            in2 => \N__1447\,
            in3 => \N__2433\,
            lcout => \uart_tx.M_bitCtr_qZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNIP5AF3_0_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2384\,
            in1 => \N__1848\,
            in2 => \N__2436\,
            in3 => \N__1920\,
            lcout => \uart_tx.N_143_0\,
            ltout => \uart_tx.N_143_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_1_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__1871\,
            in1 => \_gnd_net_\,
            in2 => \N__1444\,
            in3 => \N__2311\,
            lcout => \uart_tx.M_bitCtr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNITA5V2_0_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2426\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1918\,
            lcout => OPEN,
            ltout => \uart_tx_N_185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_RNIE6EK8_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__1522\,
            in1 => \N__2309\,
            in2 => \N__1441\,
            in3 => \N__1555\,
            lcout => OPEN,
            ltout => \click_dtct_M_count_d6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_0_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100000011"
        )
    port map (
            in0 => \N__2310\,
            in1 => \N__1483\,
            in2 => \N__1561\,
            in3 => \N__1588\,
            lcout => \uart_tx.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNITT1L_1_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__1870\,
            in1 => \N__1845\,
            in2 => \_gnd_net_\,
            in3 => \N__2425\,
            lcout => OPEN,
            ltout => \uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNIUE4P3_2_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2383\,
            in1 => \N__1804\,
            in2 => \N__1558\,
            in3 => \N__1919\,
            lcout => \uart_tx_N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_1_1_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2424\,
            in2 => \_gnd_net_\,
            in3 => \N__2382\,
            lcout => \uart_tx_N_186_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_0_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001111000"
        )
    port map (
            in0 => \N__2317\,
            in1 => \N__1585\,
            in2 => \N__2238\,
            in3 => \N__1524\,
            lcout => \M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2898\,
            ce => 'H',
            sr => \N__1497\
        );

    \M_count_q_RNITRFR_3_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2789\,
            in2 => \_gnd_net_\,
            in3 => \N__2230\,
            lcout => OPEN,
            ltout => \un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIF6FD2_1_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2818\,
            in1 => \N__2755\,
            in2 => \N__1549\,
            in3 => \N__2304\,
            lcout => \un1_M_count_q_ac0_5_m2_0_a2_3\,
            ltout => \un1_M_count_q_ac0_5_m2_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_4_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111111100000"
        )
    port map (
            in0 => \N__1587\,
            in1 => \N__1523\,
            in2 => \N__1540\,
            in3 => \N__2163\,
            lcout => \M_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2898\,
            ce => 'H',
            sr => \N__1497\
        );

    \M_count_q_1_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001111000"
        )
    port map (
            in0 => \N__1537\,
            in1 => \N__1586\,
            in2 => \N__2766\,
            in3 => \N__1525\,
            lcout => \M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2898\,
            ce => 'H',
            sr => \N__1497\
        );

    \btn_cond.M_ctr_q_RNIUMNB_4_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2664\,
            in1 => \N__2682\,
            in2 => \N__2626\,
            in3 => \N__2645\,
            lcout => \btn_cond.out_17_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNO_0_7_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__2714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2198\,
            lcout => \un1_M_count_q_axbxc7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIE6NB_0_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3096\,
            in1 => \N__3158\,
            in2 => \N__3121\,
            in3 => \N__3138\,
            lcout => btn_cond_out_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIQGM2_12_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3055\,
            in1 => \N__3072\,
            in2 => \N__2521\,
            in3 => \N__2498\,
            lcout => OPEN,
            ltout => \btn_cond.out_17_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIKBLL_10_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1567\,
            in2 => \N__1600\,
            in3 => \N__1597\,
            lcout => btn_cond_out_17,
            ltout => \btn_cond_out_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_RNIUTK51_0_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__2004\,
            in1 => \N__2062\,
            in2 => \N__1591\,
            in3 => \N__2091\,
            lcout => click_dtct_out8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__2063\,
            in1 => \_gnd_net_\,
            in2 => \N__2095\,
            in3 => \N__2032\,
            lcout => \click_dtct_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIA1N2_19_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3007\,
            in1 => \N__2984\,
            in2 => \N__2965\,
            in3 => \N__3024\,
            lcout => btn_cond_out_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIS377_10_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2602\,
            in1 => \N__2558\,
            in2 => \N__2581\,
            in3 => \N__2538\,
            lcout => \btn_cond.out_17_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_0_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1762\,
            lcout => \reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_2_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1729\,
            lcout => \reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_1_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1763\,
            in2 => \_gnd_net_\,
            in3 => \N__1735\,
            lcout => \reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_0_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2314\,
            in1 => \N__1708\,
            in2 => \N__1723\,
            in3 => \N__1722\,
            lcout => \uart_tx.M_ctr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_0\,
            clk => \N__2893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2327\,
            in1 => \N__1695\,
            in2 => \_gnd_net_\,
            in3 => \N__1681\,
            lcout => \uart_tx.M_ctr_qZ1Z_1\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_0\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_1\,
            clk => \N__2893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_2_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1678\,
            in2 => \_gnd_net_\,
            in3 => \N__1660\,
            lcout => \uart_tx.M_ctr_q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_1\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_3_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2328\,
            in1 => \N__1657\,
            in2 => \_gnd_net_\,
            in3 => \N__1645\,
            lcout => \uart_tx.M_ctr_qZ0Z_3\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_2\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_3\,
            clk => \N__2893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_4_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2315\,
            in1 => \N__1642\,
            in2 => \_gnd_net_\,
            in3 => \N__1630\,
            lcout => \uart_tx.M_ctr_qZ1Z_4\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_3\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_4\,
            clk => \N__2893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_5_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1627\,
            in2 => \_gnd_net_\,
            in3 => \N__1609\,
            lcout => \uart_tx.M_ctr_q_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_4\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_6_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1894\,
            in2 => \_gnd_net_\,
            in3 => \N__1945\,
            lcout => OPEN,
            ltout => \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_6_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__1941\,
            in1 => \N__2316\,
            in2 => \N__1927\,
            in3 => \N__1924\,
            lcout => \uart_tx.M_ctr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_2_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__1803\,
            in1 => \N__1873\,
            in2 => \N__1882\,
            in3 => \N__2323\,
            lcout => \uart_tx.M_bitCtr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_2_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2773\,
            in1 => \N__2836\,
            in2 => \_gnd_net_\,
            in3 => \N__1802\,
            lcout => \uart_tx.M_txReg_q_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_4_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__1800\,
            in1 => \N__2146\,
            in2 => \_gnd_net_\,
            in3 => \N__2212\,
            lcout => OPEN,
            ltout => \uart_tx.M_txReg_q_RNOZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_3_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__1872\,
            in1 => \N__1846\,
            in2 => \N__1855\,
            in3 => \N__1780\,
            lcout => OPEN,
            ltout => \uart_tx.M_txReg_d_3_7_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_0_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__1847\,
            in1 => \N__1822\,
            in2 => \N__1813\,
            in3 => \N__1810\,
            lcout => \uart_tx.M_txReg_d_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_1_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__1801\,
            in1 => \N__2701\,
            in2 => \_gnd_net_\,
            in3 => \N__2734\,
            lcout => \uart_tx.M_txReg_q_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_5_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2800\,
            in1 => \N__2176\,
            in2 => \_gnd_net_\,
            in3 => \N__1799\,
            lcout => \uart_tx.M_txReg_q_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNICJ341_19_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2089\,
            in1 => \N__2065\,
            in2 => \_gnd_net_\,
            in3 => \N__2030\,
            lcout => OPEN,
            ltout => \M_btn_cond_out_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_RNIJC4S1_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__2005\,
            in1 => \_gnd_net_\,
            in2 => \N__1966\,
            in3 => \N__2305\,
            lcout => \M_count_d6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_0_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3139\,
            in2 => \N__3175\,
            in3 => \N__3174\,
            lcout => \btn_cond.M_ctr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => \btn_cond.un1_M_ctr_q_cry_0\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_1_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3097\,
            in2 => \_gnd_net_\,
            in3 => \N__1963\,
            lcout => \btn_cond.M_ctr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_0\,
            carryout => \btn_cond.un1_M_ctr_q_cry_1\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_2_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3159\,
            in2 => \_gnd_net_\,
            in3 => \N__1960\,
            lcout => \btn_cond.M_ctr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_1\,
            carryout => \btn_cond.un1_M_ctr_q_cry_2\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_3_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3119\,
            in2 => \_gnd_net_\,
            in3 => \N__1957\,
            lcout => \btn_cond.M_ctr_qZ0Z_3\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_2\,
            carryout => \btn_cond.un1_M_ctr_q_cry_3\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_4_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2646\,
            in2 => \_gnd_net_\,
            in3 => \N__1954\,
            lcout => \btn_cond.M_ctr_qZ0Z_4\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_3\,
            carryout => \btn_cond.un1_M_ctr_q_cry_4\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_5_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2665\,
            in2 => \_gnd_net_\,
            in3 => \N__1951\,
            lcout => \btn_cond.M_ctr_qZ0Z_5\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_4\,
            carryout => \btn_cond.un1_M_ctr_q_cry_5\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_6_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2683\,
            in2 => \_gnd_net_\,
            in3 => \N__1948\,
            lcout => \btn_cond.M_ctr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_5\,
            carryout => \btn_cond.un1_M_ctr_q_cry_6\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_7_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2622\,
            in2 => \_gnd_net_\,
            in3 => \N__2122\,
            lcout => \btn_cond.M_ctr_qZ0Z_7\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_6\,
            carryout => \btn_cond.un1_M_ctr_q_cry_7\,
            clk => \N__2899\,
            ce => 'H',
            sr => \N__2461\
        );

    \btn_cond.M_ctr_q_8_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2580\,
            in2 => \_gnd_net_\,
            in3 => \N__2119\,
            lcout => \btn_cond.M_ctr_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => \btn_cond.un1_M_ctr_q_cry_8\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_9_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2539\,
            in2 => \_gnd_net_\,
            in3 => \N__2116\,
            lcout => \btn_cond.M_ctr_qZ0Z_9\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_8\,
            carryout => \btn_cond.un1_M_ctr_q_cry_9\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_10_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2559\,
            in2 => \_gnd_net_\,
            in3 => \N__2113\,
            lcout => \btn_cond.M_ctr_qZ0Z_10\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_9\,
            carryout => \btn_cond.un1_M_ctr_q_cry_10\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_11_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2601\,
            in2 => \_gnd_net_\,
            in3 => \N__2110\,
            lcout => \btn_cond.M_ctr_qZ0Z_11\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_10\,
            carryout => \btn_cond.un1_M_ctr_q_cry_11\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_12_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3073\,
            in2 => \_gnd_net_\,
            in3 => \N__2107\,
            lcout => \btn_cond.M_ctr_qZ0Z_12\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_11\,
            carryout => \btn_cond.un1_M_ctr_q_cry_12\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_13_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3051\,
            in2 => \_gnd_net_\,
            in3 => \N__2104\,
            lcout => \btn_cond.M_ctr_qZ0Z_13\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_12\,
            carryout => \btn_cond.un1_M_ctr_q_cry_13\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_14_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2500\,
            in2 => \_gnd_net_\,
            in3 => \N__2101\,
            lcout => \btn_cond.M_ctr_qZ0Z_14\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_13\,
            carryout => \btn_cond.un1_M_ctr_q_cry_14\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_15_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2520\,
            in2 => \_gnd_net_\,
            in3 => \N__2098\,
            lcout => \btn_cond.M_ctr_qZ0Z_15\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_14\,
            carryout => \btn_cond.un1_M_ctr_q_cry_15\,
            clk => \N__2902\,
            ce => 'H',
            sr => \N__2460\
        );

    \btn_cond.M_ctr_q_16_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2961\,
            in2 => \_gnd_net_\,
            in3 => \N__2473\,
            lcout => \btn_cond.M_ctr_qZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => \btn_cond.un1_M_ctr_q_cry_16\,
            clk => \N__2904\,
            ce => 'H',
            sr => \N__2459\
        );

    \btn_cond.M_ctr_q_17_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3006\,
            in2 => \_gnd_net_\,
            in3 => \N__2470\,
            lcout => \btn_cond.M_ctr_qZ0Z_17\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_16\,
            carryout => \btn_cond.un1_M_ctr_q_cry_17\,
            clk => \N__2904\,
            ce => 'H',
            sr => \N__2459\
        );

    \btn_cond.M_ctr_q_18_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3025\,
            in2 => \_gnd_net_\,
            in3 => \N__2467\,
            lcout => \btn_cond.M_ctr_qZ0Z_18\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_17\,
            carryout => \btn_cond.un1_M_ctr_q_cry_18\,
            clk => \N__2904\,
            ce => 'H',
            sr => \N__2459\
        );

    \btn_cond.M_ctr_q_19_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2985\,
            in2 => \_gnd_net_\,
            in3 => \N__2464\,
            lcout => \btn_cond.M_ctr_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2904\,
            ce => 'H',
            sr => \N__2459\
        );

    \uart_tx.M_txReg_q_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111000110011"
        )
    port map (
            in0 => \N__2446\,
            in1 => \N__2440\,
            in2 => \_gnd_net_\,
            in3 => \N__2389\,
            lcout => usb_tx_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2889\,
            ce => 'H',
            sr => \N__2329\
        );

    \uart_tx.M_savedData_q_0_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2242\,
            lcout => \uart_tx.M_savedData_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2891\,
            ce => \N__2695\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_6_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2203\,
            lcout => \uart_tx.M_savedData_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2891\,
            ce => \N__2695\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_4_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2170\,
            lcout => \uart_tx.M_savedData_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2891\,
            ce => \N__2695\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_7_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2140\,
            lcout => \uart_tx.M_savedData_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2891\,
            ce => \N__2695\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_2_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2827\,
            lcout => \uart_tx.M_savedData_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2894\,
            ce => \N__2694\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_3_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2794\,
            lcout => \uart_tx.M_savedData_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2894\,
            ce => \N__2694\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_1_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2767\,
            lcout => \uart_tx.M_savedData_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2894\,
            ce => \N__2694\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_5_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2728\,
            lcout => \uart_tx.M_savedData_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2894\,
            ce => \N__2694\,
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIUMNB_0_4_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__2681\,
            in1 => \N__2663\,
            in2 => \N__2647\,
            in3 => \N__2618\,
            lcout => \btn_cond.g0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIS377_0_10_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__2597\,
            in1 => \N__2576\,
            in2 => \N__2560\,
            in3 => \N__2537\,
            lcout => OPEN,
            ltout => \btn_cond.g0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIMKT9_14_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__2516\,
            in1 => \N__2499\,
            in2 => \N__2482\,
            in3 => \N__3031\,
            lcout => OPEN,
            ltout => \btn_cond.g0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNICJ341_14_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2479\,
            in1 => \N__3079\,
            in2 => \N__3178\,
            in3 => \N__2941\,
            lcout => \btn_cond.M_btn_cond_out_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIE6NB_0_0_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3160\,
            in1 => \N__3137\,
            in2 => \N__3120\,
            in3 => \N__3095\,
            lcout => \btn_cond.g0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIB6B1_12_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3071\,
            in2 => \_gnd_net_\,
            in3 => \N__3047\,
            lcout => \btn_cond.g0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIA1N2_0_19_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3023\,
            in1 => \N__3002\,
            in2 => \N__2986\,
            in3 => \N__2957\,
            lcout => \btn_cond.g0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.sync.M_pipe_q_1_LC_16_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2911\,
            lcout => \btn_cond.sync.M_sync_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.sync.M_pipe_q_0_LC_16_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \btn_cond.sync.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.sync.M_pipe_q_RNIJLM5_1_LC_16_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2848\,
            lcout => \btn_cond.sync.M_sync_out_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
