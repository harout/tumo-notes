-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Oct 28 2022 20:54:26

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    dout : out std_logic_vector(6 downto 0);
    usb_tx : out std_logic;
    usb_rx : in std_logic;
    sr_latch : out std_logic;
    sr_data : out std_logic;
    sr_clk : out std_logic;
    rst_n : in std_logic;
    last : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__4357\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2218\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2136\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2046\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2014\ : std_logic;
signal \N__2011\ : std_logic;
signal \N__2008\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1993\ : std_logic;
signal \N__1992\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1972\ : std_logic;
signal \N__1969\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1921\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1912\ : std_logic;
signal \N__1909\ : std_logic;
signal \N__1906\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1888\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1840\ : std_logic;
signal usb_rx_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal rst_n_c : std_logic;
signal \reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal sr_chain_latch_e1_i : std_logic;
signal \bfn_28_18_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_7_s1\ : std_logic;
signal \bfn_28_19_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_15_s1\ : std_logic;
signal \bfn_28_20_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_23_s1\ : std_logic;
signal \bfn_28_21_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1_THRU_CO\ : std_logic;
signal \sr_chain.latch_0_sqmuxa_cascade_\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_11\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_7_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_8\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_9\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_0\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_3\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_10\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_15\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_12\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_2\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_15_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_13\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_14\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_20\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_23\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_21\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_22\ : std_logic;
signal \sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_\ : std_logic;
signal \sr_chain.M_sr_bit_d_0_sqmuxa_cascade_\ : std_logic;
signal \sr_chain.un1_M_sr_clock_count_q_1_c2\ : std_logic;
signal \sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_2\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_3\ : std_logic;
signal \sr_chain.M_sr_is_sending_q_RNIMJKTZ0\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_1\ : std_logic;
signal \bfn_30_18_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_0\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_1\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_2\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_3\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_4\ : std_logic;
signal \sr_chain.M_main_clock_count_q_i_23\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_5\ : std_logic;
signal \sr_chain.M_main_clock_count_d8\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_0_and\ : std_logic;
signal \bfn_30_19_0_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_0\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_2_and\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_1\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_3_and\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_2\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_3\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_5_and\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_4\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_24\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_q_i_24\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_5\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_6\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_4\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_5\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_1_and\ : std_logic;
signal \sr_chain.M_sr_bit_d_4_6_ns_1_0\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_4\ : std_logic;
signal \sr_chain.M_sr_bit_d_1_sqmuxa_cascade_\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_7_0_cascade_\ : std_logic;
signal \sr_chain.M_sr_bit_q_3\ : std_logic;
signal dout_c_1 : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_16\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_19\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_17\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_18\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_4_and\ : std_logic;
signal \sr_chain.latch_0_sqmuxa\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1_THRU_CO\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_6\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1_THRU_CO\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\ : std_logic;
signal \sr_chain.M_sr_rest_cycles_qZ0Z_7\ : std_logic;
signal \N_100_g\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_3_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_4_and\ : std_logic;
signal \sr_chain.M_sr_bit_d_0_sqmuxa\ : std_logic;
signal \sr_chain.M_sr_data_buffer_qZ0Z_3\ : std_logic;
signal \sr_chain.M_main_clock_count_d_0_sqmuxa\ : std_logic;
signal \sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_1_and\ : std_logic;
signal \sr_chain.un1_M_sr_clock_count_q\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_THRU_CO\ : std_logic;
signal \M_reset_cond_out_0\ : std_logic;
signal \sr_chain.latch_0_sqmuxa_1_0_cascade_\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_0_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_5_and\ : std_logic;
signal \sr_chain.M_main_clock_count_d8_2_and\ : std_logic;
signal \sr_chain.M_sr_clock_count_qZ0Z_0\ : std_logic;
signal \sr_chain.latch_0_sqmuxa_1_0\ : std_logic;
signal \sr_chain.latch13\ : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\ : std_logic;
signal dout_c_0 : std_logic;
signal \sr_chain.un1_M_sr_rest_cycles_q_3_0\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_0\ : std_logic;
signal \bfn_32_17_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_1\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_0\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_2\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_1\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_3\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_2\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_4\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_3\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_5\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_4\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_6\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_5\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_7\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_6\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_7\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_8\ : std_logic;
signal \bfn_32_18_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_9\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_8\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_10\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_9\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_11\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_10\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_12\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_11\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_13\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_12\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_14\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_13\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_15\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_14\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_15\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_16\ : std_logic;
signal \bfn_32_19_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_17\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_16\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_18\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_17\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_19\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_18\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_20\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_19\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_21\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_20\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_22\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_21\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_23\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_22\ : std_logic;
signal \sr_chain.un1_M_main_clock_count_q_1_cry_23\ : std_logic;
signal \bfn_32_20_0_\ : std_logic;
signal \sr_chain.M_main_clock_count_qZ0Z_24\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_c_g : std_logic;
signal \sr_chain.N_36_g\ : std_logic;

signal clk_wire : std_logic;
signal dout_wire : std_logic_vector(6 downto 0);
signal last_wire : std_logic;
signal rst_n_wire : std_logic;
signal sr_clk_wire : std_logic;
signal sr_data_wire : std_logic;
signal sr_latch_wire : std_logic;
signal usb_rx_wire : std_logic;
signal usb_tx_wire : std_logic;

begin
    clk_wire <= clk;
    dout <= dout_wire;
    last <= last_wire;
    rst_n_wire <= rst_n;
    sr_clk <= sr_clk_wire;
    sr_data <= sr_data_wire;
    sr_latch <= sr_latch_wire;
    usb_rx_wire <= usb_rx;
    usb_tx <= usb_tx_wire;

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__4355\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4357\,
            DIN => \N__4356\,
            DOUT => \N__4355\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4357\,
            PADOUT => \N__4356\,
            PADIN => \N__4355\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \dout_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4346\,
            DIN => \N__4345\,
            DOUT => \N__4344\,
            PACKAGEPIN => dout_wire(0)
        );

    \dout_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4346\,
            PADOUT => \N__4345\,
            PADIN => \N__4344\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3376\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \dout_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4337\,
            DIN => \N__4336\,
            DOUT => \N__4335\,
            PACKAGEPIN => dout_wire(1)
        );

    \dout_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4337\,
            PADOUT => \N__4336\,
            PADIN => \N__4335\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2857\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \dout_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4328\,
            DIN => \N__4327\,
            DOUT => \N__4326\,
            PACKAGEPIN => dout_wire(2)
        );

    \dout_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4328\,
            PADOUT => \N__4327\,
            PADIN => \N__4326\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1879\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \dout_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4319\,
            DIN => \N__4318\,
            DOUT => \N__4317\,
            PACKAGEPIN => dout_wire(3)
        );

    \dout_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__4319\,
            PADOUT => \N__4318\,
            PADIN => \N__4317\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \dout_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4310\,
            DIN => \N__4309\,
            DOUT => \N__4308\,
            PACKAGEPIN => dout_wire(4)
        );

    \dout_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__4310\,
            PADOUT => \N__4309\,
            PADIN => \N__4308\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \dout_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4301\,
            DIN => \N__4300\,
            DOUT => \N__4299\,
            PACKAGEPIN => dout_wire(5)
        );

    \dout_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__4301\,
            PADOUT => \N__4300\,
            PADIN => \N__4299\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \dout_obuft_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4292\,
            DIN => \N__4291\,
            DOUT => \N__4290\,
            PACKAGEPIN => dout_wire(6)
        );

    \dout_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__4292\,
            PADOUT => \N__4291\,
            PADIN => \N__4290\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \last_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4283\,
            DIN => \N__4282\,
            DOUT => \N__4281\,
            PACKAGEPIN => last_wire
        );

    \last_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4283\,
            PADOUT => \N__4282\,
            PADIN => \N__4281\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4274\,
            DIN => \N__4273\,
            DOUT => \N__4272\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4274\,
            PADOUT => \N__4273\,
            PADIN => \N__4272\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \sr_clk_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4265\,
            DIN => \N__4264\,
            DOUT => \N__4263\,
            PACKAGEPIN => sr_clk_wire
        );

    \sr_clk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4265\,
            PADOUT => \N__4264\,
            PADIN => \N__4263\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \sr_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4256\,
            DIN => \N__4255\,
            DOUT => \N__4254\,
            PACKAGEPIN => sr_data_wire
        );

    \sr_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4256\,
            PADOUT => \N__4255\,
            PADIN => \N__4254\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \sr_latch_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4247\,
            DIN => \N__4246\,
            DOUT => \N__4245\,
            PACKAGEPIN => sr_latch_wire
        );

    \sr_latch_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4247\,
            PADOUT => \N__4246\,
            PADIN => \N__4245\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \usb_rx_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4238\,
            DIN => \N__4237\,
            DOUT => \N__4236\,
            PACKAGEPIN => usb_rx_wire
        );

    \usb_rx_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4238\,
            PADOUT => \N__4237\,
            PADIN => \N__4236\,
            CLOCKENABLE => 'H',
            DIN0 => usb_rx_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \usb_tx_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4229\,
            DIN => \N__4228\,
            DOUT => \N__4227\,
            PACKAGEPIN => usb_tx_wire
        );

    \usb_tx_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4229\,
            PADOUT => \N__4228\,
            PADIN => \N__4227\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1849\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__4210\,
            I => \N__4206\
        );

    \I__950\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4203\
        );

    \I__949\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4200\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4203\,
            I => \sr_chain.M_main_clock_count_qZ0Z_18\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4200\,
            I => \sr_chain.M_main_clock_count_qZ0Z_18\
        );

    \I__946\ : InMux
    port map (
            O => \N__4195\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_17\
        );

    \I__945\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4188\
        );

    \I__944\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4185\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4188\,
            I => \sr_chain.M_main_clock_count_qZ0Z_19\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4185\,
            I => \sr_chain.M_main_clock_count_qZ0Z_19\
        );

    \I__941\ : InMux
    port map (
            O => \N__4180\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_18\
        );

    \I__940\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4173\
        );

    \I__939\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4170\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4173\,
            I => \sr_chain.M_main_clock_count_qZ0Z_20\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4170\,
            I => \sr_chain.M_main_clock_count_qZ0Z_20\
        );

    \I__936\ : InMux
    port map (
            O => \N__4165\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_19\
        );

    \I__935\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4158\
        );

    \I__934\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4155\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4158\,
            I => \sr_chain.M_main_clock_count_qZ0Z_21\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4155\,
            I => \sr_chain.M_main_clock_count_qZ0Z_21\
        );

    \I__931\ : InMux
    port map (
            O => \N__4150\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_20\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__4147\,
            I => \N__4143\
        );

    \I__929\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4140\
        );

    \I__928\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4137\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4140\,
            I => \sr_chain.M_main_clock_count_qZ0Z_22\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4137\,
            I => \sr_chain.M_main_clock_count_qZ0Z_22\
        );

    \I__925\ : InMux
    port map (
            O => \N__4132\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_21\
        );

    \I__924\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4122\
        );

    \I__922\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4119\
        );

    \I__921\ : Span4Mux_h
    port map (
            O => \N__4122\,
            I => \N__4116\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4119\,
            I => \sr_chain.M_main_clock_count_qZ0Z_23\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__4116\,
            I => \sr_chain.M_main_clock_count_qZ0Z_23\
        );

    \I__918\ : InMux
    port map (
            O => \N__4111\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_22\
        );

    \I__917\ : InMux
    port map (
            O => \N__4108\,
            I => \bfn_32_20_0_\
        );

    \I__916\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4101\
        );

    \I__915\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4098\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4101\,
            I => \sr_chain.M_main_clock_count_qZ0Z_24\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4098\,
            I => \sr_chain.M_main_clock_count_qZ0Z_24\
        );

    \I__912\ : ClkMux
    port map (
            O => \N__4093\,
            I => \N__4042\
        );

    \I__911\ : ClkMux
    port map (
            O => \N__4092\,
            I => \N__4042\
        );

    \I__910\ : ClkMux
    port map (
            O => \N__4091\,
            I => \N__4042\
        );

    \I__909\ : ClkMux
    port map (
            O => \N__4090\,
            I => \N__4042\
        );

    \I__908\ : ClkMux
    port map (
            O => \N__4089\,
            I => \N__4042\
        );

    \I__907\ : ClkMux
    port map (
            O => \N__4088\,
            I => \N__4042\
        );

    \I__906\ : ClkMux
    port map (
            O => \N__4087\,
            I => \N__4042\
        );

    \I__905\ : ClkMux
    port map (
            O => \N__4086\,
            I => \N__4042\
        );

    \I__904\ : ClkMux
    port map (
            O => \N__4085\,
            I => \N__4042\
        );

    \I__903\ : ClkMux
    port map (
            O => \N__4084\,
            I => \N__4042\
        );

    \I__902\ : ClkMux
    port map (
            O => \N__4083\,
            I => \N__4042\
        );

    \I__901\ : ClkMux
    port map (
            O => \N__4082\,
            I => \N__4042\
        );

    \I__900\ : ClkMux
    port map (
            O => \N__4081\,
            I => \N__4042\
        );

    \I__899\ : ClkMux
    port map (
            O => \N__4080\,
            I => \N__4042\
        );

    \I__898\ : ClkMux
    port map (
            O => \N__4079\,
            I => \N__4042\
        );

    \I__897\ : ClkMux
    port map (
            O => \N__4078\,
            I => \N__4042\
        );

    \I__896\ : ClkMux
    port map (
            O => \N__4077\,
            I => \N__4042\
        );

    \I__895\ : GlobalMux
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__894\ : gio2CtrlBuf
    port map (
            O => \N__4039\,
            I => clk_c_g
        );

    \I__893\ : SRMux
    port map (
            O => \N__4036\,
            I => \N__4024\
        );

    \I__892\ : SRMux
    port map (
            O => \N__4035\,
            I => \N__4024\
        );

    \I__891\ : SRMux
    port map (
            O => \N__4034\,
            I => \N__4024\
        );

    \I__890\ : SRMux
    port map (
            O => \N__4033\,
            I => \N__4024\
        );

    \I__889\ : GlobalMux
    port map (
            O => \N__4024\,
            I => \N__4021\
        );

    \I__888\ : gio2CtrlBuf
    port map (
            O => \N__4021\,
            I => \sr_chain.N_36_g\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__4018\,
            I => \N__4014\
        );

    \I__886\ : InMux
    port map (
            O => \N__4017\,
            I => \N__4011\
        );

    \I__885\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4008\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__4003\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4008\,
            I => \N__4003\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__4003\,
            I => \sr_chain.M_main_clock_count_qZ0Z_10\
        );

    \I__881\ : InMux
    port map (
            O => \N__4000\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_9\
        );

    \I__880\ : InMux
    port map (
            O => \N__3997\,
            I => \N__3993\
        );

    \I__879\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3990\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__3993\,
            I => \sr_chain.M_main_clock_count_qZ0Z_11\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__3990\,
            I => \sr_chain.M_main_clock_count_qZ0Z_11\
        );

    \I__876\ : InMux
    port map (
            O => \N__3985\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_10\
        );

    \I__875\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3978\
        );

    \I__874\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3975\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__3978\,
            I => \sr_chain.M_main_clock_count_qZ0Z_12\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__3975\,
            I => \sr_chain.M_main_clock_count_qZ0Z_12\
        );

    \I__871\ : InMux
    port map (
            O => \N__3970\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_11\
        );

    \I__870\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3963\
        );

    \I__869\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3960\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__3963\,
            I => \sr_chain.M_main_clock_count_qZ0Z_13\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__3960\,
            I => \sr_chain.M_main_clock_count_qZ0Z_13\
        );

    \I__866\ : InMux
    port map (
            O => \N__3955\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_12\
        );

    \I__865\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3948\
        );

    \I__864\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3945\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__3948\,
            I => \sr_chain.M_main_clock_count_qZ0Z_14\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__3945\,
            I => \sr_chain.M_main_clock_count_qZ0Z_14\
        );

    \I__861\ : InMux
    port map (
            O => \N__3940\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_13\
        );

    \I__860\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3933\
        );

    \I__859\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3930\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__3933\,
            I => \N__3927\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__3930\,
            I => \sr_chain.M_main_clock_count_qZ0Z_15\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__3927\,
            I => \sr_chain.M_main_clock_count_qZ0Z_15\
        );

    \I__855\ : InMux
    port map (
            O => \N__3922\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_14\
        );

    \I__854\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3915\
        );

    \I__853\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3912\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__3915\,
            I => \sr_chain.M_main_clock_count_qZ0Z_16\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__3912\,
            I => \sr_chain.M_main_clock_count_qZ0Z_16\
        );

    \I__850\ : InMux
    port map (
            O => \N__3907\,
            I => \bfn_32_19_0_\
        );

    \I__849\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3900\
        );

    \I__848\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3897\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__3900\,
            I => \N__3894\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__3897\,
            I => \sr_chain.M_main_clock_count_qZ0Z_17\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__3894\,
            I => \sr_chain.M_main_clock_count_qZ0Z_17\
        );

    \I__844\ : InMux
    port map (
            O => \N__3889\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_16\
        );

    \I__843\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3882\
        );

    \I__842\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3879\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__3882\,
            I => \sr_chain.M_main_clock_count_qZ0Z_2\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__3879\,
            I => \sr_chain.M_main_clock_count_qZ0Z_2\
        );

    \I__839\ : InMux
    port map (
            O => \N__3874\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_1\
        );

    \I__838\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3867\
        );

    \I__837\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3864\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__3867\,
            I => \sr_chain.M_main_clock_count_qZ0Z_3\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__3864\,
            I => \sr_chain.M_main_clock_count_qZ0Z_3\
        );

    \I__834\ : InMux
    port map (
            O => \N__3859\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_2\
        );

    \I__833\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3852\
        );

    \I__832\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3849\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__3852\,
            I => \sr_chain.M_main_clock_count_qZ0Z_4\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__3849\,
            I => \sr_chain.M_main_clock_count_qZ0Z_4\
        );

    \I__829\ : InMux
    port map (
            O => \N__3844\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_3\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__3841\,
            I => \N__3837\
        );

    \I__827\ : InMux
    port map (
            O => \N__3840\,
            I => \N__3834\
        );

    \I__826\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3831\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__3834\,
            I => \sr_chain.M_main_clock_count_qZ0Z_5\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__3831\,
            I => \sr_chain.M_main_clock_count_qZ0Z_5\
        );

    \I__823\ : InMux
    port map (
            O => \N__3826\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_4\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__3823\,
            I => \N__3819\
        );

    \I__821\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3816\
        );

    \I__820\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3813\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__3816\,
            I => \sr_chain.M_main_clock_count_qZ0Z_6\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__3813\,
            I => \sr_chain.M_main_clock_count_qZ0Z_6\
        );

    \I__817\ : InMux
    port map (
            O => \N__3808\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_5\
        );

    \I__816\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3801\
        );

    \I__815\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3798\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__3801\,
            I => \N__3795\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3798\,
            I => \sr_chain.M_main_clock_count_qZ0Z_7\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__3795\,
            I => \sr_chain.M_main_clock_count_qZ0Z_7\
        );

    \I__811\ : InMux
    port map (
            O => \N__3790\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_6\
        );

    \I__810\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3783\
        );

    \I__809\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3780\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__3783\,
            I => \sr_chain.M_main_clock_count_qZ0Z_8\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__3780\,
            I => \sr_chain.M_main_clock_count_qZ0Z_8\
        );

    \I__806\ : InMux
    port map (
            O => \N__3775\,
            I => \bfn_32_18_0_\
        );

    \I__805\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3768\
        );

    \I__804\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3765\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__3768\,
            I => \sr_chain.M_main_clock_count_qZ0Z_9\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__3765\,
            I => \sr_chain.M_main_clock_count_qZ0Z_9\
        );

    \I__801\ : InMux
    port map (
            O => \N__3760\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_8\
        );

    \I__800\ : InMux
    port map (
            O => \N__3757\,
            I => \N__3752\
        );

    \I__799\ : InMux
    port map (
            O => \N__3756\,
            I => \N__3749\
        );

    \I__798\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3746\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__3752\,
            I => \N__3743\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__3749\,
            I => \sr_chain.un1_M_sr_clock_count_q\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__3746\,
            I => \sr_chain.un1_M_sr_clock_count_q\
        );

    \I__794\ : Odrv12
    port map (
            O => \N__3743\,
            I => \sr_chain.un1_M_sr_clock_count_q\
        );

    \I__793\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3732\
        );

    \I__792\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3727\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__3732\,
            I => \N__3724\
        );

    \I__790\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3721\
        );

    \I__789\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3718\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__3727\,
            I => \sr_chain.M_main_clock_count_d8_THRU_CO\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__3724\,
            I => \sr_chain.M_main_clock_count_d8_THRU_CO\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__3721\,
            I => \sr_chain.M_main_clock_count_d8_THRU_CO\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3718\,
            I => \sr_chain.M_main_clock_count_d8_THRU_CO\
        );

    \I__784\ : IoInMux
    port map (
            O => \N__3709\,
            I => \N__3704\
        );

    \I__783\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3700\
        );

    \I__782\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3697\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3704\,
            I => \N__3694\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__3703\,
            I => \N__3691\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3700\,
            I => \N__3686\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3697\,
            I => \N__3683\
        );

    \I__777\ : Span4Mux_s3_v
    port map (
            O => \N__3694\,
            I => \N__3680\
        );

    \I__776\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3671\
        );

    \I__775\ : InMux
    port map (
            O => \N__3690\,
            I => \N__3671\
        );

    \I__774\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3671\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__3686\,
            I => \N__3668\
        );

    \I__772\ : Span4Mux_v
    port map (
            O => \N__3683\,
            I => \N__3665\
        );

    \I__771\ : Sp12to4
    port map (
            O => \N__3680\,
            I => \N__3662\
        );

    \I__770\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3657\
        );

    \I__769\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3657\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3671\,
            I => \N__3654\
        );

    \I__767\ : Span4Mux_h
    port map (
            O => \N__3668\,
            I => \N__3651\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__3665\,
            I => \N__3648\
        );

    \I__765\ : Span12Mux_h
    port map (
            O => \N__3662\,
            I => \N__3645\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3657\,
            I => \N__3640\
        );

    \I__763\ : Sp12to4
    port map (
            O => \N__3654\,
            I => \N__3640\
        );

    \I__762\ : Sp12to4
    port map (
            O => \N__3651\,
            I => \N__3631\
        );

    \I__761\ : Sp12to4
    port map (
            O => \N__3648\,
            I => \N__3631\
        );

    \I__760\ : Span12Mux_v
    port map (
            O => \N__3645\,
            I => \N__3631\
        );

    \I__759\ : Span12Mux_s6_h
    port map (
            O => \N__3640\,
            I => \N__3631\
        );

    \I__758\ : Odrv12
    port map (
            O => \N__3631\,
            I => \M_reset_cond_out_0\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__3628\,
            I => \sr_chain.latch_0_sqmuxa_1_0_cascade_\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__3625\,
            I => \N__3622\
        );

    \I__755\ : InMux
    port map (
            O => \N__3622\,
            I => \N__3619\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3619\,
            I => \sr_chain.M_main_clock_count_d8_0_and\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__752\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3610\,
            I => \sr_chain.M_main_clock_count_d8_5_and\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__3607\,
            I => \N__3604\
        );

    \I__749\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__3601\,
            I => \sr_chain.M_main_clock_count_d8_2_and\
        );

    \I__747\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3592\
        );

    \I__746\ : InMux
    port map (
            O => \N__3597\,
            I => \N__3588\
        );

    \I__745\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3583\
        );

    \I__744\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3583\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3592\,
            I => \N__3580\
        );

    \I__742\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3575\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3588\,
            I => \N__3568\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3583\,
            I => \N__3568\
        );

    \I__739\ : Span4Mux_h
    port map (
            O => \N__3580\,
            I => \N__3568\
        );

    \I__738\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3563\
        );

    \I__737\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3563\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3575\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_0\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3568\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_0\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3563\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_0\
        );

    \I__733\ : InMux
    port map (
            O => \N__3556\,
            I => \N__3553\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3553\,
            I => \sr_chain.latch_0_sqmuxa_1_0\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__3550\,
            I => \N__3544\
        );

    \I__730\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3538\
        );

    \I__729\ : InMux
    port map (
            O => \N__3548\,
            I => \N__3538\
        );

    \I__728\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3534\
        );

    \I__727\ : InMux
    port map (
            O => \N__3544\,
            I => \N__3529\
        );

    \I__726\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3526\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3538\,
            I => \N__3523\
        );

    \I__724\ : InMux
    port map (
            O => \N__3537\,
            I => \N__3520\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3534\,
            I => \N__3517\
        );

    \I__722\ : InMux
    port map (
            O => \N__3533\,
            I => \N__3514\
        );

    \I__721\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3511\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__3529\,
            I => \sr_chain.latch13\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3526\,
            I => \sr_chain.latch13\
        );

    \I__718\ : Odrv4
    port map (
            O => \N__3523\,
            I => \sr_chain.latch13\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3520\,
            I => \sr_chain.latch13\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__3517\,
            I => \sr_chain.latch13\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3514\,
            I => \sr_chain.latch13\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3511\,
            I => \sr_chain.latch13\
        );

    \I__713\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3483\
        );

    \I__712\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3479\
        );

    \I__711\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3474\
        );

    \I__710\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3474\
        );

    \I__709\ : InMux
    port map (
            O => \N__3492\,
            I => \N__3471\
        );

    \I__708\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3461\
        );

    \I__707\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3458\
        );

    \I__706\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3449\
        );

    \I__705\ : InMux
    port map (
            O => \N__3488\,
            I => \N__3449\
        );

    \I__704\ : InMux
    port map (
            O => \N__3487\,
            I => \N__3449\
        );

    \I__703\ : InMux
    port map (
            O => \N__3486\,
            I => \N__3449\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3483\,
            I => \N__3446\
        );

    \I__701\ : InMux
    port map (
            O => \N__3482\,
            I => \N__3443\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3479\,
            I => \N__3438\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3474\,
            I => \N__3438\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3471\,
            I => \N__3435\
        );

    \I__697\ : InMux
    port map (
            O => \N__3470\,
            I => \N__3430\
        );

    \I__696\ : InMux
    port map (
            O => \N__3469\,
            I => \N__3427\
        );

    \I__695\ : InMux
    port map (
            O => \N__3468\,
            I => \N__3424\
        );

    \I__694\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3415\
        );

    \I__693\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3415\
        );

    \I__692\ : InMux
    port map (
            O => \N__3465\,
            I => \N__3415\
        );

    \I__691\ : InMux
    port map (
            O => \N__3464\,
            I => \N__3415\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3461\,
            I => \N__3406\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3458\,
            I => \N__3406\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3449\,
            I => \N__3406\
        );

    \I__687\ : Span4Mux_h
    port map (
            O => \N__3446\,
            I => \N__3406\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3443\,
            I => \N__3403\
        );

    \I__685\ : Span4Mux_h
    port map (
            O => \N__3438\,
            I => \N__3398\
        );

    \I__684\ : Span4Mux_s1_h
    port map (
            O => \N__3435\,
            I => \N__3398\
        );

    \I__683\ : InMux
    port map (
            O => \N__3434\,
            I => \N__3393\
        );

    \I__682\ : InMux
    port map (
            O => \N__3433\,
            I => \N__3393\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3430\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3427\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3424\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3415\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__3406\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__3403\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__3398\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3393\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\
        );

    \I__673\ : IoInMux
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__671\ : IoSpan4Mux
    port map (
            O => \N__3370\,
            I => \N__3367\
        );

    \I__670\ : Span4Mux_s1_h
    port map (
            O => \N__3367\,
            I => \N__3364\
        );

    \I__669\ : Sp12to4
    port map (
            O => \N__3364\,
            I => \N__3361\
        );

    \I__668\ : Span12Mux_s9_h
    port map (
            O => \N__3361\,
            I => \N__3358\
        );

    \I__667\ : Span12Mux_h
    port map (
            O => \N__3358\,
            I => \N__3355\
        );

    \I__666\ : Odrv12
    port map (
            O => \N__3355\,
            I => dout_c_0
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__3352\,
            I => \N__3348\
        );

    \I__664\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3345\
        );

    \I__663\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3342\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3345\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_3_0\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3342\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_3_0\
        );

    \I__660\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3333\
        );

    \I__659\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3330\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3333\,
            I => \sr_chain.M_main_clock_count_qZ0Z_0\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3330\,
            I => \sr_chain.M_main_clock_count_qZ0Z_0\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__3325\,
            I => \N__3321\
        );

    \I__655\ : InMux
    port map (
            O => \N__3324\,
            I => \N__3318\
        );

    \I__654\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3315\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3318\,
            I => \sr_chain.M_main_clock_count_qZ0Z_1\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3315\,
            I => \sr_chain.M_main_clock_count_qZ0Z_1\
        );

    \I__651\ : InMux
    port map (
            O => \N__3310\,
            I => \sr_chain.un1_M_main_clock_count_q_1_cry_0\
        );

    \I__650\ : InMux
    port map (
            O => \N__3307\,
            I => \N__3301\
        );

    \I__649\ : InMux
    port map (
            O => \N__3306\,
            I => \N__3298\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__3305\,
            I => \N__3295\
        );

    \I__647\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3285\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3301\,
            I => \N__3280\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3298\,
            I => \N__3280\
        );

    \I__644\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3271\
        );

    \I__643\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3271\
        );

    \I__642\ : InMux
    port map (
            O => \N__3293\,
            I => \N__3271\
        );

    \I__641\ : InMux
    port map (
            O => \N__3292\,
            I => \N__3271\
        );

    \I__640\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3262\
        );

    \I__639\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3262\
        );

    \I__638\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3262\
        );

    \I__637\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3262\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3285\,
            I => \N__3252\
        );

    \I__635\ : Span4Mux_h
    port map (
            O => \N__3280\,
            I => \N__3252\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3271\,
            I => \N__3252\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3262\,
            I => \N__3252\
        );

    \I__632\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3249\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3252\,
            I => \sr_chain.latch_0_sqmuxa\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3249\,
            I => \sr_chain.latch_0_sqmuxa\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__628\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3238\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3238\,
            I => \N__3235\
        );

    \I__626\ : Span4Mux_s3_h
    port map (
            O => \N__3235\,
            I => \N__3232\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__3232\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1_THRU_CO\
        );

    \I__624\ : InMux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3226\,
            I => \N__3222\
        );

    \I__622\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3218\
        );

    \I__621\ : Span4Mux_h
    port map (
            O => \N__3222\,
            I => \N__3215\
        );

    \I__620\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3212\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3218\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_6\
        );

    \I__618\ : Odrv4
    port map (
            O => \N__3215\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_6\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3212\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_6\
        );

    \I__616\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3202\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__614\ : Span4Mux_s3_h
    port map (
            O => \N__3199\,
            I => \N__3196\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__3196\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1_THRU_CO\
        );

    \I__612\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3182\
        );

    \I__611\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3182\
        );

    \I__610\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3173\
        );

    \I__609\ : InMux
    port map (
            O => \N__3190\,
            I => \N__3173\
        );

    \I__608\ : InMux
    port map (
            O => \N__3189\,
            I => \N__3173\
        );

    \I__607\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3173\
        );

    \I__606\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3166\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3182\,
            I => \N__3162\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3173\,
            I => \N__3159\
        );

    \I__603\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3150\
        );

    \I__602\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3150\
        );

    \I__601\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3150\
        );

    \I__600\ : InMux
    port map (
            O => \N__3169\,
            I => \N__3150\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3166\,
            I => \N__3147\
        );

    \I__598\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3144\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__3162\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__3159\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3150\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__594\ : Odrv4
    port map (
            O => \N__3147\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3144\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\
        );

    \I__592\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3130\,
            I => \N__3126\
        );

    \I__590\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3122\
        );

    \I__589\ : Span4Mux_h
    port map (
            O => \N__3126\,
            I => \N__3119\
        );

    \I__588\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3116\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3122\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_7\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__3119\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_7\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3116\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_7\
        );

    \I__584\ : SRMux
    port map (
            O => \N__3109\,
            I => \N__3088\
        );

    \I__583\ : SRMux
    port map (
            O => \N__3108\,
            I => \N__3088\
        );

    \I__582\ : SRMux
    port map (
            O => \N__3107\,
            I => \N__3088\
        );

    \I__581\ : SRMux
    port map (
            O => \N__3106\,
            I => \N__3088\
        );

    \I__580\ : SRMux
    port map (
            O => \N__3105\,
            I => \N__3088\
        );

    \I__579\ : SRMux
    port map (
            O => \N__3104\,
            I => \N__3088\
        );

    \I__578\ : SRMux
    port map (
            O => \N__3103\,
            I => \N__3088\
        );

    \I__577\ : GlobalMux
    port map (
            O => \N__3088\,
            I => \N__3085\
        );

    \I__576\ : gio2CtrlBuf
    port map (
            O => \N__3085\,
            I => \N_100_g\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__574\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3076\,
            I => \sr_chain.M_main_clock_count_d8_3_and\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__3073\,
            I => \N__3070\
        );

    \I__571\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3067\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3067\,
            I => \sr_chain.M_main_clock_count_d8_4_and\
        );

    \I__569\ : InMux
    port map (
            O => \N__3064\,
            I => \N__3059\
        );

    \I__568\ : InMux
    port map (
            O => \N__3063\,
            I => \N__3054\
        );

    \I__567\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3054\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3059\,
            I => \sr_chain.M_sr_bit_d_0_sqmuxa\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3054\,
            I => \sr_chain.M_sr_bit_d_0_sqmuxa\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3049\,
            I => \N__3046\
        );

    \I__563\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3042\
        );

    \I__562\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3039\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3042\,
            I => \N__3036\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3039\,
            I => \N__3031\
        );

    \I__559\ : Span4Mux_h
    port map (
            O => \N__3036\,
            I => \N__3031\
        );

    \I__558\ : Odrv4
    port map (
            O => \N__3031\,
            I => \sr_chain.M_sr_data_buffer_qZ0Z_3\
        );

    \I__557\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3023\
        );

    \I__556\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3018\
        );

    \I__555\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3018\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3023\,
            I => \sr_chain.M_main_clock_count_d_0_sqmuxa\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3018\,
            I => \sr_chain.M_main_clock_count_d_0_sqmuxa\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__3013\,
            I => \sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_\
        );

    \I__551\ : IoInMux
    port map (
            O => \N__3010\,
            I => \N__3007\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3007\,
            I => \N__3004\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__3004\,
            I => \sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3001\,
            I => \N__2998\
        );

    \I__547\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2995\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2995\,
            I => \sr_chain.M_main_clock_count_d8_1_and\
        );

    \I__545\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2988\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__2991\,
            I => \N__2985\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2988\,
            I => \N__2982\
        );

    \I__542\ : InMux
    port map (
            O => \N__2985\,
            I => \N__2979\
        );

    \I__541\ : Span4Mux_s3_h
    port map (
            O => \N__2982\,
            I => \N__2976\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2979\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_24\
        );

    \I__539\ : Odrv4
    port map (
            O => \N__2976\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_24\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__2971\,
            I => \N__2968\
        );

    \I__537\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2965\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2965\,
            I => \sr_chain.M_sr_rest_cycles_q_i_24\
        );

    \I__535\ : InMux
    port map (
            O => \N__2962\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_6\
        );

    \I__534\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2955\
        );

    \I__533\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2951\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2955\,
            I => \N__2948\
        );

    \I__531\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2945\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__2951\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_4\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__2948\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_4\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__2945\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_4\
        );

    \I__527\ : InMux
    port map (
            O => \N__2938\,
            I => \N__2933\
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__2937\,
            I => \N__2930\
        );

    \I__525\ : InMux
    port map (
            O => \N__2936\,
            I => \N__2927\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__2933\,
            I => \N__2924\
        );

    \I__523\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2921\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2927\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_5\
        );

    \I__521\ : Odrv4
    port map (
            O => \N__2924\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_5\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__2921\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_5\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__2914\,
            I => \N__2911\
        );

    \I__518\ : InMux
    port map (
            O => \N__2911\,
            I => \N__2908\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__2908\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_1_and\
        );

    \I__516\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2902\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__2902\,
            I => \N__2899\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__2899\,
            I => \sr_chain.M_sr_bit_d_4_6_ns_1_0\
        );

    \I__513\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2892\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__2895\,
            I => \N__2889\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__2892\,
            I => \N__2886\
        );

    \I__510\ : InMux
    port map (
            O => \N__2889\,
            I => \N__2882\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__2886\,
            I => \N__2879\
        );

    \I__508\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2876\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__2882\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_4\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__2879\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_4\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__2876\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_4\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__2869\,
            I => \sr_chain.M_sr_bit_d_1_sqmuxa_cascade_\
        );

    \I__503\ : CascadeMux
    port map (
            O => \N__2866\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_7_0_cascade_\
        );

    \I__502\ : InMux
    port map (
            O => \N__2863\,
            I => \N__2860\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2860\,
            I => \sr_chain.M_sr_bit_q_3\
        );

    \I__500\ : IoInMux
    port map (
            O => \N__2857\,
            I => \N__2854\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2854\,
            I => \N__2851\
        );

    \I__498\ : Span12Mux_s8_h
    port map (
            O => \N__2851\,
            I => \N__2848\
        );

    \I__497\ : Span12Mux_h
    port map (
            O => \N__2848\,
            I => \N__2844\
        );

    \I__496\ : InMux
    port map (
            O => \N__2847\,
            I => \N__2841\
        );

    \I__495\ : Odrv12
    port map (
            O => \N__2844\,
            I => dout_c_1
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2841\,
            I => dout_c_1
        );

    \I__493\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2831\
        );

    \I__492\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2828\
        );

    \I__491\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2825\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2831\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_16\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2828\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_16\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__2825\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_16\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__2818\,
            I => \N__2815\
        );

    \I__486\ : InMux
    port map (
            O => \N__2815\,
            I => \N__2810\
        );

    \I__485\ : InMux
    port map (
            O => \N__2814\,
            I => \N__2807\
        );

    \I__484\ : InMux
    port map (
            O => \N__2813\,
            I => \N__2804\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2810\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_19\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__2807\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_19\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2804\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_19\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__2797\,
            I => \N__2792\
        );

    \I__479\ : InMux
    port map (
            O => \N__2796\,
            I => \N__2789\
        );

    \I__478\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2786\
        );

    \I__477\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2783\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2789\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_17\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2786\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_17\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2783\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_17\
        );

    \I__473\ : CascadeMux
    port map (
            O => \N__2776\,
            I => \N__2773\
        );

    \I__472\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2768\
        );

    \I__471\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2765\
        );

    \I__470\ : InMux
    port map (
            O => \N__2771\,
            I => \N__2762\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2768\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_18\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2765\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_18\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2762\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_18\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__2755\,
            I => \N__2752\
        );

    \I__465\ : InMux
    port map (
            O => \N__2752\,
            I => \N__2749\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2749\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_4_and\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__2746\,
            I => \N__2743\
        );

    \I__462\ : InMux
    port map (
            O => \N__2743\,
            I => \N__2740\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__2740\,
            I => \sr_chain.M_main_clock_count_q_i_23\
        );

    \I__460\ : InMux
    port map (
            O => \N__2737\,
            I => \sr_chain.M_main_clock_count_d8\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__458\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2728\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_0_and\
        );

    \I__456\ : CascadeMux
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__455\ : InMux
    port map (
            O => \N__2722\,
            I => \N__2719\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2719\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_2_and\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__2716\,
            I => \N__2713\
        );

    \I__452\ : InMux
    port map (
            O => \N__2713\,
            I => \N__2710\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2710\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_3_and\
        );

    \I__450\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2704\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2704\,
            I => \N__2701\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__2701\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_1_5_and\
        );

    \I__447\ : InMux
    port map (
            O => \N__2698\,
            I => \N__2692\
        );

    \I__446\ : InMux
    port map (
            O => \N__2697\,
            I => \N__2692\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2692\,
            I => \sr_chain.un1_M_sr_clock_count_q_1_c2\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__2689\,
            I => \sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_\
        );

    \I__443\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2679\
        );

    \I__442\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2674\
        );

    \I__441\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2674\
        );

    \I__440\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2669\
        );

    \I__439\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2669\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2679\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_2\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2674\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_2\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2669\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_2\
        );

    \I__435\ : InMux
    port map (
            O => \N__2662\,
            I => \N__2654\
        );

    \I__434\ : InMux
    port map (
            O => \N__2661\,
            I => \N__2654\
        );

    \I__433\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2649\
        );

    \I__432\ : InMux
    port map (
            O => \N__2659\,
            I => \N__2649\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2654\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_3\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2649\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_3\
        );

    \I__429\ : SRMux
    port map (
            O => \N__2644\,
            I => \N__2641\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2641\,
            I => \N__2637\
        );

    \I__427\ : InMux
    port map (
            O => \N__2640\,
            I => \N__2634\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__2637\,
            I => \sr_chain.M_sr_is_sending_q_RNIMJKTZ0\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2634\,
            I => \sr_chain.M_sr_is_sending_q_RNIMJKTZ0\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__2629\,
            I => \N__2625\
        );

    \I__423\ : CascadeMux
    port map (
            O => \N__2628\,
            I => \N__2622\
        );

    \I__422\ : InMux
    port map (
            O => \N__2625\,
            I => \N__2617\
        );

    \I__421\ : InMux
    port map (
            O => \N__2622\,
            I => \N__2610\
        );

    \I__420\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2610\
        );

    \I__419\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2610\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2617\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_1\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2610\,
            I => \sr_chain.M_sr_clock_count_qZ0Z_1\
        );

    \I__416\ : InMux
    port map (
            O => \N__2605\,
            I => \N__2602\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2602\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1_THRU_CO\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__413\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2593\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2593\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1_THRU_CO\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__2590\,
            I => \N__2587\
        );

    \I__410\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2582\
        );

    \I__409\ : InMux
    port map (
            O => \N__2586\,
            I => \N__2577\
        );

    \I__408\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2577\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2582\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_20\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2577\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_20\
        );

    \I__405\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2567\
        );

    \I__404\ : InMux
    port map (
            O => \N__2571\,
            I => \N__2564\
        );

    \I__403\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2561\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2567\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_23\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2564\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_23\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2561\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_23\
        );

    \I__399\ : CascadeMux
    port map (
            O => \N__2554\,
            I => \N__2551\
        );

    \I__398\ : InMux
    port map (
            O => \N__2551\,
            I => \N__2548\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2548\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1_THRU_CO\
        );

    \I__396\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2540\
        );

    \I__395\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2537\
        );

    \I__394\ : InMux
    port map (
            O => \N__2543\,
            I => \N__2534\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2540\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_21\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2537\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_21\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2534\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_21\
        );

    \I__390\ : InMux
    port map (
            O => \N__2527\,
            I => \N__2524\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2524\,
            I => \N__2521\
        );

    \I__388\ : Odrv4
    port map (
            O => \N__2521\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1_THRU_CO\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__2518\,
            I => \N__2513\
        );

    \I__386\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2510\
        );

    \I__385\ : InMux
    port map (
            O => \N__2516\,
            I => \N__2507\
        );

    \I__384\ : InMux
    port map (
            O => \N__2513\,
            I => \N__2504\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2510\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_22\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2507\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_22\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2504\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_22\
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__2497\,
            I => \sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__2494\,
            I => \sr_chain.M_sr_bit_d_0_sqmuxa_cascade_\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__2491\,
            I => \N__2488\
        );

    \I__377\ : InMux
    port map (
            O => \N__2488\,
            I => \N__2485\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2485\,
            I => \N__2482\
        );

    \I__375\ : Odrv4
    port map (
            O => \N__2482\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1_THRU_CO\
        );

    \I__374\ : InMux
    port map (
            O => \N__2479\,
            I => \N__2474\
        );

    \I__373\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2469\
        );

    \I__372\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2469\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2474\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_12\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2469\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_12\
        );

    \I__369\ : InMux
    port map (
            O => \N__2464\,
            I => \N__2461\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2461\,
            I => \N__2458\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__2458\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1_THRU_CO\
        );

    \I__366\ : InMux
    port map (
            O => \N__2455\,
            I => \N__2451\
        );

    \I__365\ : InMux
    port map (
            O => \N__2454\,
            I => \N__2447\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2451\,
            I => \N__2444\
        );

    \I__363\ : InMux
    port map (
            O => \N__2450\,
            I => \N__2441\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2447\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_2\
        );

    \I__361\ : Odrv4
    port map (
            O => \N__2444\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_2\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2441\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_2\
        );

    \I__359\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2431\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2431\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1_THRU_CO\
        );

    \I__357\ : InMux
    port map (
            O => \N__2428\,
            I => \N__2425\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2425\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1_THRU_CO\
        );

    \I__355\ : InMux
    port map (
            O => \N__2422\,
            I => \N__2419\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2419\,
            I => \N__2416\
        );

    \I__353\ : Odrv4
    port map (
            O => \N__2416\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1_THRU_CO\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__2413\,
            I => \N__2410\
        );

    \I__351\ : InMux
    port map (
            O => \N__2410\,
            I => \N__2407\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2407\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_15_s1_THRU_CO\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__2404\,
            I => \N__2401\
        );

    \I__348\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2398\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2398\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1_THRU_CO\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__2395\,
            I => \N__2390\
        );

    \I__345\ : InMux
    port map (
            O => \N__2394\,
            I => \N__2387\
        );

    \I__344\ : InMux
    port map (
            O => \N__2393\,
            I => \N__2384\
        );

    \I__343\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2381\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2387\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_13\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2384\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_13\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2381\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_13\
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__2374\,
            I => \N__2371\
        );

    \I__338\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2368\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2368\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1_THRU_CO\
        );

    \I__336\ : InMux
    port map (
            O => \N__2365\,
            I => \N__2360\
        );

    \I__335\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2357\
        );

    \I__334\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2354\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2360\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_14\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2357\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_14\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2354\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_14\
        );

    \I__330\ : InMux
    port map (
            O => \N__2347\,
            I => \N__2344\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2344\,
            I => \N__2341\
        );

    \I__328\ : Span4Mux_h
    port map (
            O => \N__2341\,
            I => \N__2338\
        );

    \I__327\ : Odrv4
    port map (
            O => \N__2338\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1_THRU_CO\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2335\,
            I => \N__2332\
        );

    \I__325\ : InMux
    port map (
            O => \N__2332\,
            I => \N__2329\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2329\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_7_s1_THRU_CO\
        );

    \I__323\ : InMux
    port map (
            O => \N__2326\,
            I => \N__2321\
        );

    \I__322\ : InMux
    port map (
            O => \N__2325\,
            I => \N__2316\
        );

    \I__321\ : InMux
    port map (
            O => \N__2324\,
            I => \N__2316\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2321\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_8\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2316\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_8\
        );

    \I__318\ : InMux
    port map (
            O => \N__2311\,
            I => \N__2308\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2308\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1_THRU_CO\
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__2305\,
            I => \N__2301\
        );

    \I__315\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2297\
        );

    \I__314\ : InMux
    port map (
            O => \N__2301\,
            I => \N__2292\
        );

    \I__313\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2292\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2297\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_9\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2292\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_9\
        );

    \I__310\ : InMux
    port map (
            O => \N__2287\,
            I => \N__2283\
        );

    \I__309\ : InMux
    port map (
            O => \N__2286\,
            I => \N__2280\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2283\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_0\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2280\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_0\
        );

    \I__306\ : InMux
    port map (
            O => \N__2275\,
            I => \N__2272\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2272\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1_THRU_CO\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2269\,
            I => \N__2264\
        );

    \I__303\ : InMux
    port map (
            O => \N__2268\,
            I => \N__2261\
        );

    \I__302\ : InMux
    port map (
            O => \N__2267\,
            I => \N__2258\
        );

    \I__301\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2255\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2261\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_1\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2258\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_1\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2255\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_1\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__2248\,
            I => \N__2245\
        );

    \I__296\ : InMux
    port map (
            O => \N__2245\,
            I => \N__2242\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2242\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1_THRU_CO\
        );

    \I__294\ : InMux
    port map (
            O => \N__2239\,
            I => \N__2234\
        );

    \I__293\ : InMux
    port map (
            O => \N__2238\,
            I => \N__2231\
        );

    \I__292\ : InMux
    port map (
            O => \N__2237\,
            I => \N__2228\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2234\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_3\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2231\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_3\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2228\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_3\
        );

    \I__288\ : InMux
    port map (
            O => \N__2221\,
            I => \N__2218\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2218\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1_THRU_CO\
        );

    \I__286\ : InMux
    port map (
            O => \N__2215\,
            I => \N__2210\
        );

    \I__285\ : InMux
    port map (
            O => \N__2214\,
            I => \N__2207\
        );

    \I__284\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2204\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2210\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_10\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2207\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_10\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2204\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_10\
        );

    \I__280\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2194\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2194\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1_THRU_CO\
        );

    \I__278\ : CascadeMux
    port map (
            O => \N__2191\,
            I => \N__2188\
        );

    \I__277\ : InMux
    port map (
            O => \N__2188\,
            I => \N__2183\
        );

    \I__276\ : InMux
    port map (
            O => \N__2187\,
            I => \N__2178\
        );

    \I__275\ : InMux
    port map (
            O => \N__2186\,
            I => \N__2178\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2183\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_15\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2178\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_15\
        );

    \I__272\ : InMux
    port map (
            O => \N__2173\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1\
        );

    \I__271\ : CascadeMux
    port map (
            O => \N__2170\,
            I => \N__2161\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__2169\,
            I => \N__2158\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__2168\,
            I => \N__2155\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__2167\,
            I => \N__2152\
        );

    \I__267\ : CascadeMux
    port map (
            O => \N__2166\,
            I => \N__2149\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__2165\,
            I => \N__2146\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__2164\,
            I => \N__2143\
        );

    \I__264\ : InMux
    port map (
            O => \N__2161\,
            I => \N__2129\
        );

    \I__263\ : InMux
    port map (
            O => \N__2158\,
            I => \N__2129\
        );

    \I__262\ : InMux
    port map (
            O => \N__2155\,
            I => \N__2129\
        );

    \I__261\ : InMux
    port map (
            O => \N__2152\,
            I => \N__2120\
        );

    \I__260\ : InMux
    port map (
            O => \N__2149\,
            I => \N__2120\
        );

    \I__259\ : InMux
    port map (
            O => \N__2146\,
            I => \N__2120\
        );

    \I__258\ : InMux
    port map (
            O => \N__2143\,
            I => \N__2120\
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__2142\,
            I => \N__2117\
        );

    \I__256\ : CascadeMux
    port map (
            O => \N__2141\,
            I => \N__2114\
        );

    \I__255\ : CascadeMux
    port map (
            O => \N__2140\,
            I => \N__2111\
        );

    \I__254\ : CascadeMux
    port map (
            O => \N__2139\,
            I => \N__2101\
        );

    \I__253\ : CascadeMux
    port map (
            O => \N__2138\,
            I => \N__2098\
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__2137\,
            I => \N__2094\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__2136\,
            I => \N__2091\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2129\,
            I => \N__2086\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2120\,
            I => \N__2086\
        );

    \I__248\ : InMux
    port map (
            O => \N__2117\,
            I => \N__2079\
        );

    \I__247\ : InMux
    port map (
            O => \N__2114\,
            I => \N__2079\
        );

    \I__246\ : InMux
    port map (
            O => \N__2111\,
            I => \N__2079\
        );

    \I__245\ : CascadeMux
    port map (
            O => \N__2110\,
            I => \N__2076\
        );

    \I__244\ : CascadeMux
    port map (
            O => \N__2109\,
            I => \N__2073\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2108\,
            I => \N__2069\
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__2107\,
            I => \N__2066\
        );

    \I__241\ : CascadeMux
    port map (
            O => \N__2106\,
            I => \N__2063\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__2105\,
            I => \N__2060\
        );

    \I__239\ : CascadeMux
    port map (
            O => \N__2104\,
            I => \N__2057\
        );

    \I__238\ : InMux
    port map (
            O => \N__2101\,
            I => \N__2046\
        );

    \I__237\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2046\
        );

    \I__236\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2046\
        );

    \I__235\ : InMux
    port map (
            O => \N__2094\,
            I => \N__2046\
        );

    \I__234\ : InMux
    port map (
            O => \N__2091\,
            I => \N__2046\
        );

    \I__233\ : Span4Mux_h
    port map (
            O => \N__2086\,
            I => \N__2041\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2079\,
            I => \N__2041\
        );

    \I__231\ : InMux
    port map (
            O => \N__2076\,
            I => \N__2030\
        );

    \I__230\ : InMux
    port map (
            O => \N__2073\,
            I => \N__2030\
        );

    \I__229\ : InMux
    port map (
            O => \N__2072\,
            I => \N__2030\
        );

    \I__228\ : InMux
    port map (
            O => \N__2069\,
            I => \N__2030\
        );

    \I__227\ : InMux
    port map (
            O => \N__2066\,
            I => \N__2030\
        );

    \I__226\ : InMux
    port map (
            O => \N__2063\,
            I => \N__2023\
        );

    \I__225\ : InMux
    port map (
            O => \N__2060\,
            I => \N__2023\
        );

    \I__224\ : InMux
    port map (
            O => \N__2057\,
            I => \N__2023\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2046\,
            I => \CONSTANT_ONE_NET\
        );

    \I__222\ : Odrv4
    port map (
            O => \N__2041\,
            I => \CONSTANT_ONE_NET\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2030\,
            I => \CONSTANT_ONE_NET\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2023\,
            I => \CONSTANT_ONE_NET\
        );

    \I__219\ : InMux
    port map (
            O => \N__2014\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1\
        );

    \I__218\ : InMux
    port map (
            O => \N__2011\,
            I => \bfn_28_21_0_\
        );

    \I__217\ : InMux
    port map (
            O => \N__2008\,
            I => \N__2005\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__2005\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1_THRU_CO\
        );

    \I__215\ : InMux
    port map (
            O => \N__2002\,
            I => \N__1999\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1999\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1_THRU_CO\
        );

    \I__213\ : CascadeMux
    port map (
            O => \N__1996\,
            I => \sr_chain.latch_0_sqmuxa_cascade_\
        );

    \I__212\ : CascadeMux
    port map (
            O => \N__1993\,
            I => \N__1988\
        );

    \I__211\ : InMux
    port map (
            O => \N__1992\,
            I => \N__1985\
        );

    \I__210\ : InMux
    port map (
            O => \N__1991\,
            I => \N__1982\
        );

    \I__209\ : InMux
    port map (
            O => \N__1988\,
            I => \N__1979\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1985\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_11\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1982\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_11\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1979\,
            I => \sr_chain.M_sr_rest_cycles_qZ0Z_11\
        );

    \I__205\ : InMux
    port map (
            O => \N__1972\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1\
        );

    \I__204\ : InMux
    port map (
            O => \N__1969\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1\
        );

    \I__203\ : InMux
    port map (
            O => \N__1966\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1\
        );

    \I__202\ : InMux
    port map (
            O => \N__1963\,
            I => \bfn_28_20_0_\
        );

    \I__201\ : InMux
    port map (
            O => \N__1960\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1\
        );

    \I__200\ : InMux
    port map (
            O => \N__1957\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1\
        );

    \I__199\ : InMux
    port map (
            O => \N__1954\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1\
        );

    \I__198\ : InMux
    port map (
            O => \N__1951\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1\
        );

    \I__197\ : InMux
    port map (
            O => \N__1948\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1\
        );

    \I__196\ : InMux
    port map (
            O => \N__1945\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1\
        );

    \I__195\ : InMux
    port map (
            O => \N__1942\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1\
        );

    \I__194\ : InMux
    port map (
            O => \N__1939\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1\
        );

    \I__193\ : InMux
    port map (
            O => \N__1936\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1\
        );

    \I__192\ : InMux
    port map (
            O => \N__1933\,
            I => \bfn_28_19_0_\
        );

    \I__191\ : InMux
    port map (
            O => \N__1930\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1\
        );

    \I__190\ : InMux
    port map (
            O => \N__1927\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1\
        );

    \I__189\ : InMux
    port map (
            O => \N__1924\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1\
        );

    \I__188\ : InMux
    port map (
            O => \N__1921\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1\
        );

    \I__187\ : InMux
    port map (
            O => \N__1918\,
            I => \N__1915\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1915\,
            I => \reset_cond.M_stage_qZ0Z_1\
        );

    \I__185\ : InMux
    port map (
            O => \N__1912\,
            I => \N__1909\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1909\,
            I => \reset_cond.M_stage_qZ0Z_0\
        );

    \I__183\ : InMux
    port map (
            O => \N__1906\,
            I => \N__1894\
        );

    \I__182\ : InMux
    port map (
            O => \N__1905\,
            I => \N__1894\
        );

    \I__181\ : InMux
    port map (
            O => \N__1904\,
            I => \N__1894\
        );

    \I__180\ : InMux
    port map (
            O => \N__1903\,
            I => \N__1894\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1894\,
            I => \N__1891\
        );

    \I__178\ : Span12Mux_v
    port map (
            O => \N__1891\,
            I => \N__1888\
        );

    \I__177\ : Odrv12
    port map (
            O => \N__1888\,
            I => rst_n_c
        );

    \I__176\ : InMux
    port map (
            O => \N__1885\,
            I => \N__1882\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1882\,
            I => \reset_cond.M_stage_qZ0Z_2\
        );

    \I__174\ : IoInMux
    port map (
            O => \N__1879\,
            I => \N__1876\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1876\,
            I => \N__1873\
        );

    \I__172\ : Span4Mux_s3_h
    port map (
            O => \N__1873\,
            I => \N__1870\
        );

    \I__171\ : Span4Mux_v
    port map (
            O => \N__1870\,
            I => \N__1867\
        );

    \I__170\ : Sp12to4
    port map (
            O => \N__1867\,
            I => \N__1864\
        );

    \I__169\ : Span12Mux_h
    port map (
            O => \N__1864\,
            I => \N__1861\
        );

    \I__168\ : Odrv12
    port map (
            O => \N__1861\,
            I => sr_chain_latch_e1_i
        );

    \I__167\ : InMux
    port map (
            O => \N__1858\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1\
        );

    \I__166\ : InMux
    port map (
            O => \N__1855\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1\
        );

    \I__165\ : InMux
    port map (
            O => \N__1852\,
            I => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1\
        );

    \I__164\ : IoInMux
    port map (
            O => \N__1849\,
            I => \N__1846\
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1846\,
            I => \N__1843\
        );

    \I__162\ : Span12Mux_s0_v
    port map (
            O => \N__1843\,
            I => \N__1840\
        );

    \I__161\ : Odrv12
    port map (
            O => \N__1840\,
            I => usb_rx_c
        );

    \IN_MUX_bfv_30_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_30_19_0_\
        );

    \IN_MUX_bfv_30_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_30_18_0_\
        );

    \IN_MUX_bfv_28_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_28_18_0_\
        );

    \IN_MUX_bfv_28_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_7_s1\,
            carryinitout => \bfn_28_19_0_\
        );

    \IN_MUX_bfv_28_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_15_s1\,
            carryinitout => \bfn_28_20_0_\
        );

    \IN_MUX_bfv_28_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_23_s1\,
            carryinitout => \bfn_28_21_0_\
        );

    \IN_MUX_bfv_32_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_32_17_0_\
        );

    \IN_MUX_bfv_32_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_main_clock_count_q_1_cry_7\,
            carryinitout => \bfn_32_18_0_\
        );

    \IN_MUX_bfv_32_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_main_clock_count_q_1_cry_15\,
            carryinitout => \bfn_32_19_0_\
        );

    \IN_MUX_bfv_32_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sr_chain.un1_M_main_clock_count_q_1_cry_23\,
            carryinitout => \bfn_32_20_0_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3010\,
            GLOBALBUFFEROUTPUT => \sr_chain.N_36_g\
        );

    \reset_cond.M_stage_q_RNIFG9D_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3709\,
            GLOBALBUFFEROUTPUT => \N_100_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \reset_cond.M_stage_q_1_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1904\,
            in2 => \_gnd_net_\,
            in3 => \N__1912\,
            lcout => \reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_2_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1905\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1918\,
            lcout => \reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_0_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1903\,
            lcout => \reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_3_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1906\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1885\,
            lcout => \M_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_27_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIH9O82_LC_27_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3307\,
            in2 => \_gnd_net_\,
            in3 => \N__3495\,
            lcout => sr_chain_latch_e1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_0_LC_28_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2287\,
            in2 => \_gnd_net_\,
            in3 => \N__3496\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_28_18_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1\,
            clk => \N__4078\,
            ce => 'H',
            sr => \N__3107\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1_THRU_LUT4_0_LC_28_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2267\,
            in2 => \N__2164\,
            in3 => \N__1858\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_0_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1_THRU_LUT4_0_LC_28_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2455\,
            in2 => \N__2168\,
            in3 => \N__1855\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_1_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1_THRU_LUT4_0_LC_28_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2238\,
            in2 => \N__2165\,
            in3 => \N__1852\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_2_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1_THRU_LUT4_0_LC_28_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2959\,
            in2 => \N__2169\,
            in3 => \N__1945\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_3_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1_THRU_LUT4_0_LC_28_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2938\,
            in2 => \N__2166\,
            in3 => \N__1942\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_4_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1_THRU_LUT4_0_LC_28_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3229\,
            in2 => \N__2170\,
            in3 => \N__1939\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_5_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1_THRU_LUT4_0_LC_28_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3133\,
            in2 => \N__2167\,
            in3 => \N__1936\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_6_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_7_s1_THRU_LUT4_0_LC_28_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2326\,
            in2 => \N__2138\,
            in3 => \N__1933\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_7_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_28_19_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1_THRU_LUT4_0_LC_28_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2304\,
            in2 => \N__2142\,
            in3 => \N__1930\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_8_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1_THRU_LUT4_0_LC_28_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2214\,
            in2 => \N__2139\,
            in3 => \N__1927\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_9_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1_THRU_LUT4_0_LC_28_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1991\,
            in2 => \N__2140\,
            in3 => \N__1924\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_10_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1_THRU_LUT4_0_LC_28_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2479\,
            in2 => \N__2136\,
            in3 => \N__1921\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_11_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1_THRU_LUT4_0_LC_28_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2393\,
            in2 => \N__2141\,
            in3 => \N__1972\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_12_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1_THRU_LUT4_0_LC_28_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2364\,
            in2 => \N__2137\,
            in3 => \N__1969\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_13_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1_THRU_LUT4_0_LC_28_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2097\,
            in2 => \N__2191\,
            in3 => \N__1966\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_14_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_15_s1_THRU_LUT4_0_LC_28_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2835\,
            in2 => \N__2104\,
            in3 => \N__1963\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_15_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_28_20_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1_THRU_LUT4_0_LC_28_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2795\,
            in2 => \N__2107\,
            in3 => \N__1960\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_16_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1_THRU_LUT4_0_LC_28_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2772\,
            in2 => \N__2105\,
            in3 => \N__1957\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_17_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1_THRU_LUT4_0_LC_28_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2814\,
            in2 => \N__2108\,
            in3 => \N__1954\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_18_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1_THRU_LUT4_0_LC_28_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2072\,
            in2 => \N__2590\,
            in3 => \N__1951\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_19_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1_THRU_LUT4_0_LC_28_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2544\,
            in2 => \N__2109\,
            in3 => \N__1948\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_20_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1_THRU_LUT4_0_LC_28_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2516\,
            in2 => \N__2106\,
            in3 => \N__2173\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_21_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1_THRU_LUT4_0_LC_28_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2571\,
            in2 => \N__2110\,
            in3 => \N__2014\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_22_s1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_9_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_24_LC_28_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011001011"
        )
    port map (
            in0 => \N__3306\,
            in1 => \N__3494\,
            in2 => \N__2991\,
            in3 => \N__2011\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4084\,
            ce => 'H',
            sr => \N__3103\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_RNIFAS5_LC_28_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3493\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_6_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_23_LC_28_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__2008\,
            in1 => \N__3165\,
            in2 => \_gnd_net_\,
            in3 => \N__2572\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4084\,
            ce => 'H',
            sr => \N__3103\
        );

    \sr_chain.M_sr_clock_count_q_4_LC_29_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__2685\,
            in1 => \N__2662\,
            in2 => \N__2895\,
            in3 => \N__2698\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4079\,
            ce => 'H',
            sr => \N__2644\
        );

    \sr_chain.M_sr_clock_count_q_3_LC_29_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2684\,
            in1 => \N__2661\,
            in2 => \_gnd_net_\,
            in3 => \N__2697\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4079\,
            ce => 'H',
            sr => \N__2644\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNI2VR22_LC_29_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__3755\,
            in1 => \N__3547\,
            in2 => \_gnd_net_\,
            in3 => \N__3731\,
            lcout => \sr_chain.latch_0_sqmuxa\,
            ltout => \sr_chain.latch_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_11_LC_29_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010011001"
        )
    port map (
            in0 => \N__1992\,
            in1 => \N__2002\,
            in2 => \N__1996\,
            in3 => \N__3469\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4080\,
            ce => 'H',
            sr => \N__3109\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_RNO_LC_29_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2300\,
            in1 => \N__2213\,
            in2 => \N__1993\,
            in3 => \N__2324\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_8_LC_29_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010110101010"
        )
    port map (
            in0 => \N__2325\,
            in1 => \_gnd_net_\,
            in2 => \N__2335\,
            in3 => \N__3192\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4080\,
            ce => 'H',
            sr => \N__3109\
        );

    \sr_chain.M_sr_rest_cycles_q_9_LC_29_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001011010010"
        )
    port map (
            in0 => \N__3193\,
            in1 => \N__2311\,
            in2 => \N__2305\,
            in3 => \_gnd_net_\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4080\,
            ce => 'H',
            sr => \N__3109\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_RNO_LC_29_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2237\,
            in1 => \N__2286\,
            in2 => \N__2269\,
            in3 => \N__2450\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_1_LC_29_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__2268\,
            in1 => \N__2275\,
            in2 => \_gnd_net_\,
            in3 => \N__3190\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4082\,
            ce => 'H',
            sr => \N__3108\
        );

    \sr_chain.M_sr_rest_cycles_q_3_LC_29_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010110101010"
        )
    port map (
            in0 => \N__2239\,
            in1 => \_gnd_net_\,
            in2 => \N__2248\,
            in3 => \N__3191\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4082\,
            ce => 'H',
            sr => \N__3108\
        );

    \sr_chain.M_sr_rest_cycles_q_10_LC_29_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__3188\,
            in1 => \N__2221\,
            in2 => \_gnd_net_\,
            in3 => \N__2215\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4082\,
            ce => 'H',
            sr => \N__3108\
        );

    \sr_chain.M_sr_rest_cycles_q_15_LC_29_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__2187\,
            in1 => \N__2197\,
            in2 => \_gnd_net_\,
            in3 => \N__3189\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4082\,
            ce => 'H',
            sr => \N__3108\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_RNO_LC_29_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2363\,
            in1 => \N__2186\,
            in2 => \N__2395\,
            in3 => \N__2477\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_12_LC_29_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010100101"
        )
    port map (
            in0 => \N__2478\,
            in1 => \N__3261\,
            in2 => \N__2491\,
            in3 => \N__3468\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4082\,
            ce => 'H',
            sr => \N__3108\
        );

    \sr_chain.M_sr_rest_cycles_q_2_LC_29_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__3170\,
            in1 => \N__2464\,
            in2 => \_gnd_net_\,
            in3 => \N__2454\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_17_LC_29_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__2434\,
            in1 => \N__3169\,
            in2 => \_gnd_net_\,
            in3 => \N__2796\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_19_LC_29_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010101101"
        )
    port map (
            in0 => \N__3466\,
            in1 => \N__3291\,
            in2 => \N__2818\,
            in3 => \N__2428\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_4_LC_29_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__2958\,
            in1 => \N__3171\,
            in2 => \_gnd_net_\,
            in3 => \N__2422\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_16_LC_29_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010001101"
        )
    port map (
            in0 => \N__3465\,
            in1 => \N__3290\,
            in2 => \N__2413\,
            in3 => \N__2836\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_13_LC_29_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__3288\,
            in1 => \N__2394\,
            in2 => \N__2404\,
            in3 => \N__3467\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_14_LC_29_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010001101"
        )
    port map (
            in0 => \N__3464\,
            in1 => \N__3289\,
            in2 => \N__2374\,
            in3 => \N__2365\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_5_LC_29_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__2347\,
            in1 => \N__3172\,
            in2 => \_gnd_net_\,
            in3 => \N__2936\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4085\,
            ce => 'H',
            sr => \N__3105\
        );

    \sr_chain.M_sr_rest_cycles_q_18_LC_29_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010100101"
        )
    port map (
            in0 => \N__2605\,
            in1 => \N__3292\,
            in2 => \N__2776\,
            in3 => \N__3487\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4088\,
            ce => 'H',
            sr => \N__3104\
        );

    \sr_chain.M_sr_rest_cycles_q_20_LC_29_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010100101"
        )
    port map (
            in0 => \N__2586\,
            in1 => \N__3293\,
            in2 => \N__2599\,
            in3 => \N__3488\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4088\,
            ce => 'H',
            sr => \N__3104\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_RNO_LC_29_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2543\,
            in1 => \N__2585\,
            in2 => \N__2518\,
            in3 => \N__2570\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_21_LC_29_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010100101"
        )
    port map (
            in0 => \N__2545\,
            in1 => \N__3294\,
            in2 => \N__2554\,
            in3 => \N__3489\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4088\,
            ce => 'H',
            sr => \N__3104\
        );

    \sr_chain.M_sr_rest_cycles_q_22_LC_29_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010110001"
        )
    port map (
            in0 => \N__3486\,
            in1 => \N__2527\,
            in2 => \N__3305\,
            in3 => \N__2517\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4088\,
            ce => 'H',
            sr => \N__3104\
        );

    \sr_chain.M_sr_clock_count_q_RNI63IL_1_LC_30_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2659\,
            in2 => \_gnd_net_\,
            in3 => \N__2620\,
            lcout => OPEN,
            ltout => \sr_chain.un1_M_sr_clock_count_qlto3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_RNIV7TL1_4_LC_30_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__3578\,
            in1 => \N__2885\,
            in2 => \N__2497\,
            in3 => \N__2682\,
            lcout => \sr_chain.un1_M_sr_clock_count_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_is_sending_q_RNI73BG_0_LC_30_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3537\,
            in2 => \_gnd_net_\,
            in3 => \N__3482\,
            lcout => \sr_chain.M_sr_bit_d_0_sqmuxa\,
            ltout => \sr_chain.M_sr_bit_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_is_sending_q_RNIMJKT_LC_30_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2494\,
            in3 => \N__3678\,
            lcout => \sr_chain.M_sr_is_sending_q_RNIMJKTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_RNIL1D81_1_LC_30_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3595\,
            in1 => \N__2621\,
            in2 => \_gnd_net_\,
            in3 => \N__3026\,
            lcout => \sr_chain.un1_M_sr_clock_count_q_1_c2\,
            ltout => \sr_chain.un1_M_sr_clock_count_q_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_2_LC_30_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__2686\,
            in1 => \N__3679\,
            in2 => \N__2689\,
            in3 => \N__3064\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_bit_q_RNO_2_LC_30_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111011000"
        )
    port map (
            in0 => \N__2683\,
            in1 => \N__2660\,
            in2 => \N__2629\,
            in3 => \N__3579\,
            lcout => \sr_chain.M_sr_bit_d_4_6_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_1_LC_30_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__3027\,
            in1 => \N__3596\,
            in2 => \N__2628\,
            in3 => \N__2640\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_0_c_LC_30_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3625\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_30_18_0_\,
            carryout => \sr_chain.M_main_clock_count_d8_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_1_c_LC_30_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3001\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_0\,
            carryout => \sr_chain.M_main_clock_count_d8_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_2_c_LC_30_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3607\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_1\,
            carryout => \sr_chain.M_main_clock_count_d8_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_3_c_LC_30_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_2\,
            carryout => \sr_chain.M_main_clock_count_d8_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_4_c_LC_30_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3073\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_3\,
            carryout => \sr_chain.M_main_clock_count_d8_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_5_c_LC_30_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3616\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_4\,
            carryout => \sr_chain.M_main_clock_count_d8_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_inv_LC_30_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2746\,
            in3 => \N__4129\,
            lcout => \sr_chain.M_main_clock_count_q_i_23\,
            ltout => OPEN,
            carryin => \sr_chain.M_main_clock_count_d8_5\,
            carryout => \sr_chain.M_main_clock_count_d8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_THRU_LUT4_0_LC_30_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2737\,
            lcout => \sr_chain.M_main_clock_count_d8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_0_c_LC_30_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2734\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_30_19_0_\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_LC_30_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2914\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_0\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_2_c_LC_30_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2725\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_1\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_3_c_LC_30_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2716\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_2\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_LC_30_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2755\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_3\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_5_c_LC_30_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2707\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_4\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_6_c_inv_LC_30_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2971\,
            in3 => \N__2992\,
            lcout => \sr_chain.M_sr_rest_cycles_q_i_24\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_sr_rest_cycles_q_1_5\,
            carryout => \sr_chain.un1_M_sr_rest_cycles_q_1_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_LUT4_0_LC_30_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2962\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_1_c_RNO_LC_30_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2954\,
            in1 => \N__3125\,
            in2 => \N__2937\,
            in3 => \N__3221\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_bit_q_RNO_0_LC_30_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111010"
        )
    port map (
            in0 => \N__3548\,
            in1 => \N__2905\,
            in2 => \N__3049\,
            in3 => \N__3757\,
            lcout => \sr_chain.M_sr_bit_q_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_bit_q_RNO_3_LC_30_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2896\,
            in2 => \_gnd_net_\,
            in3 => \N__3598\,
            lcout => OPEN,
            ltout => \sr_chain.M_sr_bit_d_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_bit_q_RNO_1_LC_30_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__3549\,
            in1 => \N__3736\,
            in2 => \N__2869\,
            in3 => \N__3490\,
            lcout => OPEN,
            ltout => \sr_chain.un1_M_sr_rest_cycles_q_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_bit_q_LC_30_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__2847\,
            in1 => \N__3708\,
            in2 => \N__2866\,
            in3 => \N__2863\,
            lcout => dout_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.un1_M_sr_rest_cycles_q_1_4_c_RNO_LC_30_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2834\,
            in1 => \N__2813\,
            in2 => \N__2797\,
            in3 => \N__2771\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_1_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_rest_cycles_q_6_LC_30_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000011"
        )
    port map (
            in0 => \N__3304\,
            in1 => \N__3225\,
            in2 => \N__3244\,
            in3 => \N__3491\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4091\,
            ce => 'H',
            sr => \N__3106\
        );

    \sr_chain.M_sr_rest_cycles_q_7_LC_30_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__3205\,
            in1 => \N__3187\,
            in2 => \_gnd_net_\,
            in3 => \N__3129\,
            lcout => \sr_chain.M_sr_rest_cycles_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4091\,
            ce => 'H',
            sr => \N__3106\
        );

    \sr_chain.M_main_clock_count_d8_3_c_RNO_LC_31_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3885\,
            in1 => \N__3870\,
            in2 => \N__3325\,
            in3 => \N__3336\,
            lcout => \sr_chain.M_main_clock_count_d8_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_4_c_RNO_LC_31_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3805\,
            in1 => \N__3786\,
            in2 => \N__3841\,
            in3 => \N__3855\,
            lcout => \sr_chain.M_main_clock_count_d8_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_0_LC_31_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__3063\,
            in1 => \N__3591\,
            in2 => \N__3703\,
            in3 => \N__3028\,
            lcout => \sr_chain.M_sr_clock_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_data_buffer_q_3_LC_31_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__3045\,
            in1 => \N__3690\,
            in2 => \_gnd_net_\,
            in3 => \N__3062\,
            lcout => \sr_chain.M_sr_data_buffer_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNII1RI_LC_31_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__3492\,
            in1 => \N__3533\,
            in2 => \_gnd_net_\,
            in3 => \N__3730\,
            lcout => \sr_chain.M_main_clock_count_d_0_sqmuxa\,
            ltout => \sr_chain.M_main_clock_count_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNI1I401_LC_31_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3013\,
            in3 => \N__3689\,
            lcout => \sr_chain.M_main_clock_count_d8_6_c_RNI1IZ0Z401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_1_c_RNO_LC_31_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3918\,
            in1 => \N__3951\,
            in2 => \N__4210\,
            in3 => \N__4191\,
            lcout => \sr_chain.M_main_clock_count_d8_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_6_c_RNIA6DO1_LC_31_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3756\,
            in2 => \_gnd_net_\,
            in3 => \N__3735\,
            lcout => \sr_chain.latch_0_sqmuxa_1_0\,
            ltout => \sr_chain.latch_0_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_is_sending_q_LC_31_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100010"
        )
    port map (
            in0 => \N__3434\,
            in1 => \N__3707\,
            in2 => \N__3628\,
            in3 => \N__3543\,
            lcout => \sr_chain.latch13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_0_c_RNO_LC_31_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3981\,
            in1 => \N__3966\,
            in2 => \N__3823\,
            in3 => \N__3996\,
            lcout => \sr_chain.M_main_clock_count_d8_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_is_sending_q_RNI73BG_LC_31_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3532\,
            in2 => \_gnd_net_\,
            in3 => \N__3433\,
            lcout => \sr_chain.un1_M_sr_rest_cycles_q_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_5_c_RNO_LC_31_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3937\,
            in1 => \N__3904\,
            in2 => \N__4018\,
            in3 => \N__3771\,
            lcout => \sr_chain.M_main_clock_count_d8_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_d8_2_c_RNO_LC_31_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4176\,
            in1 => \N__4104\,
            in2 => \N__4147\,
            in3 => \N__4161\,
            lcout => \sr_chain.M_main_clock_count_d8_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_sr_clock_count_q_RNI29HJ2_0_LC_31_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__3597\,
            in1 => \N__3556\,
            in2 => \N__3550\,
            in3 => \N__3470\,
            lcout => dout_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sr_chain.M_main_clock_count_q_0_LC_32_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3337\,
            in2 => \N__3352\,
            in3 => \N__3351\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_32_17_0_\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_0\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_1_LC_32_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3324\,
            in2 => \_gnd_net_\,
            in3 => \N__3310\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_0\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_1\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_2_LC_32_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3886\,
            in2 => \_gnd_net_\,
            in3 => \N__3874\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_1\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_2\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_3_LC_32_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3871\,
            in2 => \_gnd_net_\,
            in3 => \N__3859\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_2\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_3\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_4_LC_32_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3856\,
            in2 => \_gnd_net_\,
            in3 => \N__3844\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_3\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_4\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_5_LC_32_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3840\,
            in2 => \_gnd_net_\,
            in3 => \N__3826\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_4\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_5\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_6_LC_32_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3822\,
            in2 => \_gnd_net_\,
            in3 => \N__3808\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_5\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_6\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_7_LC_32_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3804\,
            in2 => \_gnd_net_\,
            in3 => \N__3790\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_6\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_7\,
            clk => \N__4087\,
            ce => 'H',
            sr => \N__4033\
        );

    \sr_chain.M_main_clock_count_q_8_LC_32_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3787\,
            in2 => \_gnd_net_\,
            in3 => \N__3775\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_32_18_0_\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_8\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_9_LC_32_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3772\,
            in2 => \_gnd_net_\,
            in3 => \N__3760\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_8\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_9\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_10_LC_32_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4017\,
            in2 => \_gnd_net_\,
            in3 => \N__4000\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_9\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_10\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_11_LC_32_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3997\,
            in2 => \_gnd_net_\,
            in3 => \N__3985\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_10\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_11\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_12_LC_32_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3982\,
            in2 => \_gnd_net_\,
            in3 => \N__3970\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_11\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_12\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_13_LC_32_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3967\,
            in2 => \_gnd_net_\,
            in3 => \N__3955\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_12\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_13\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_14_LC_32_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3952\,
            in2 => \_gnd_net_\,
            in3 => \N__3940\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_14\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_13\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_14\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_15_LC_32_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3936\,
            in2 => \_gnd_net_\,
            in3 => \N__3922\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_15\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_14\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_15\,
            clk => \N__4090\,
            ce => 'H',
            sr => \N__4034\
        );

    \sr_chain.M_main_clock_count_q_16_LC_32_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3919\,
            in2 => \_gnd_net_\,
            in3 => \N__3907\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_32_19_0_\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_16\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_17_LC_32_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3903\,
            in2 => \_gnd_net_\,
            in3 => \N__3889\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_17\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_16\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_17\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_18_LC_32_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4209\,
            in2 => \_gnd_net_\,
            in3 => \N__4195\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_18\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_17\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_18\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_19_LC_32_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4192\,
            in2 => \_gnd_net_\,
            in3 => \N__4180\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_19\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_18\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_19\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_20_LC_32_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4177\,
            in2 => \_gnd_net_\,
            in3 => \N__4165\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_20\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_19\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_20\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_21_LC_32_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4162\,
            in2 => \_gnd_net_\,
            in3 => \N__4150\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_21\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_20\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_21\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_22_LC_32_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4146\,
            in2 => \_gnd_net_\,
            in3 => \N__4132\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_22\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_21\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_22\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_23_LC_32_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4125\,
            in2 => \_gnd_net_\,
            in3 => \N__4111\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_23\,
            ltout => OPEN,
            carryin => \sr_chain.un1_M_main_clock_count_q_1_cry_22\,
            carryout => \sr_chain.un1_M_main_clock_count_q_1_cry_23\,
            clk => \N__4092\,
            ce => 'H',
            sr => \N__4035\
        );

    \sr_chain.M_main_clock_count_q_24_LC_32_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4105\,
            in2 => \_gnd_net_\,
            in3 => \N__4108\,
            lcout => \sr_chain.M_main_clock_count_qZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4093\,
            ce => 'H',
            sr => \N__4036\
        );
end \INTERFACE\;
