-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Oct 30 2022 13:51:57

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    led : out std_logic_vector(7 downto 0);
    usb_tx : out std_logic;
    trigger : in std_logic;
    rst_n : in std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__3479\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2123\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2015\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1981\ : std_logic;
signal \N__1978\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1972\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1952\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1947\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1921\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1889\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1883\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1875\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1862\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1857\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1830\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1815\ : std_logic;
signal \N__1812\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1796\ : std_logic;
signal \N__1795\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1792\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1784\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1772\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1766\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1760\ : std_logic;
signal \N__1757\ : std_logic;
signal \N__1754\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1748\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1744\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1736\ : std_logic;
signal \N__1735\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1694\ : std_logic;
signal \N__1691\ : std_logic;
signal \N__1688\ : std_logic;
signal \N__1685\ : std_logic;
signal \N__1684\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1658\ : std_logic;
signal \N__1657\ : std_logic;
signal \N__1654\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1637\ : std_logic;
signal \N__1636\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1630\ : std_logic;
signal \N__1625\ : std_logic;
signal \N__1622\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1613\ : std_logic;
signal \N__1610\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1604\ : std_logic;
signal \N__1601\ : std_logic;
signal \N__1598\ : std_logic;
signal \N__1595\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1591\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1576\ : std_logic;
signal \N__1573\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1565\ : std_logic;
signal \N__1562\ : std_logic;
signal \N__1559\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1538\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1534\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1524\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1481\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1475\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1436\ : std_logic;
signal \N__1433\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1394\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal usb_tx_c : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_4_cascade_\ : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_5\ : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_2\ : std_logic;
signal \uart_tx.M_txReg_d_3_7_ns_1_cascade_\ : std_logic;
signal \uart_tx.M_txReg_q_RNOZ0Z_1\ : std_logic;
signal \uart_tx.M_txReg_d_3\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_5\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_2\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_0\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_3\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_1\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_4\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_6\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_7\ : std_logic;
signal led_c_7 : std_logic;
signal \un1_M_count_q_axbxc7_1\ : std_logic;
signal trigger_c : std_logic;
signal \btn_cond.sync.M_sync_out_i_0\ : std_logic;
signal \btn_cond.sync.M_pipe_qZ0Z_0\ : std_logic;
signal \btn_cond.sync.M_sync_out_0\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_0\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_1\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_2\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_3\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_4\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_5\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_0\ : std_logic;
signal \uart_tx.M_ctr_qZ1Z_1\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_6\ : std_logic;
signal \uart_tx.M_ctr_qZ1Z_4\ : std_logic;
signal \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_3\ : std_logic;
signal \uart_tx.N_182_0_cascade_\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_2\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_2\ : std_logic;
signal \uart_tx.N_143_0\ : std_logic;
signal \uart_tx.N_143_0_cascade_\ : std_logic;
signal \uart_tx.N_134_i\ : std_logic;
signal \uart_tx.N_134_i_cascade_\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_5\ : std_logic;
signal \uart_tx.M_ctr_qZ1Z_5\ : std_logic;
signal \M_btn_cond_out_0_cascade_\ : std_logic;
signal \M_count_d6\ : std_logic;
signal \uart_tx.M_bitCtr_qZ0Z_1\ : std_logic;
signal \uart_tx.M_bitCtr_qZ0Z_2\ : std_logic;
signal \uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_\ : std_logic;
signal \uart_tx.N_182_0\ : std_logic;
signal \uart_tx.M_bitCtr_qZ1Z_0\ : std_logic;
signal \uart_tx_N_185\ : std_logic;
signal \click_dtct_out3_cascade_\ : std_logic;
signal \uart_tx_N_187\ : std_logic;
signal \un1_M_count_q_ac0_1\ : std_logic;
signal \un1_M_count_q_ac0_1_cascade_\ : std_logic;
signal \un1_M_count_q_ac0_7\ : std_logic;
signal \un1_M_count_q_ac0_7_cascade_\ : std_logic;
signal led_c_5 : std_logic;
signal led_c_6 : std_logic;
signal \btn_cond_out_16_5_cascade_\ : std_logic;
signal click_dtct_out_d : std_logic;
signal \btn_cond.out_17_8_cascade_\ : std_logic;
signal \btn_cond.out_17_6\ : std_logic;
signal \btn_cond.out_17_7\ : std_logic;
signal \btn_cond.g0_13_cascade_\ : std_logic;
signal \btn_cond.g0_5\ : std_logic;
signal \btn_cond.g0_14\ : std_logic;
signal \btn_cond.g0_11\ : std_logic;
signal \btn_cond.g0_16_cascade_\ : std_logic;
signal \btn_cond.g0_10\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal rst_n_c : std_logic;
signal \reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \uart_tx.N_186_1_i\ : std_logic;
signal \click_dtct_M_count_d6_0_1\ : std_logic;
signal \uart_tx.M_state_qZ0Z_1\ : std_logic;
signal \uart_tx.M_state_qZ0Z_0\ : std_logic;
signal \uart_tx_N_186_1_cascade_\ : std_logic;
signal \un1_M_count_q_ac0_out\ : std_logic;
signal led_c_3 : std_logic;
signal led_c_2 : std_logic;
signal \un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_\ : std_logic;
signal led_c_1 : std_logic;
signal \un1_M_count_q_ac0_5_m2_0_a2_3\ : std_logic;
signal \un1_M_count_q_ac0_5_m2_0_a2_3_cascade_\ : std_logic;
signal led_c_4 : std_logic;
signal btn_cond_out_16_5 : std_logic;
signal btn_cond_out_16_4 : std_logic;
signal \click_dtct_M_last_q\ : std_logic;
signal btn_cond_out_17 : std_logic;
signal click_dtct_out8 : std_logic;
signal click_dtct_out3 : std_logic;
signal \click_dtct_out8_cascade_\ : std_logic;
signal \uart_tx_N_186_1\ : std_logic;
signal led_c_0 : std_logic;
signal \M_reset_cond_out_0\ : std_logic;
signal \btn_cond.M_btn_cond_out_i_0\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_0\ : std_logic;
signal \bfn_18_27_0_\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_1\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_0\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_2\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_1\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_3\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_2\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_4\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_3\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_5\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_4\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_6\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_5\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_7\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_6\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_7\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_8\ : std_logic;
signal \bfn_18_28_0_\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_9\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_8\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_10\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_9\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_11\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_10\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_12\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_11\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_13\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_12\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_14\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_13\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_15\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_14\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_15\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_16\ : std_logic;
signal \bfn_18_29_0_\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_17\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_16\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_18\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_17\ : std_logic;
signal \btn_cond.un1_M_ctr_q_cry_18\ : std_logic;
signal \btn_cond.M_ctr_qZ0Z_19\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_c_g : std_logic;
signal \btn_cond.M_sync_out_i_g_0\ : std_logic;

signal clk_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal rst_n_wire : std_logic;
signal trigger_wire : std_logic;
signal usb_tx_wire : std_logic;

begin
    clk_wire <= clk;
    led <= led_wire;
    rst_n_wire <= rst_n;
    trigger_wire <= trigger;
    usb_tx <= usb_tx_wire;

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3477\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3479\,
            DIN => \N__3478\,
            DOUT => \N__3477\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3479\,
            PADOUT => \N__3478\,
            PADIN => \N__3477\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3468\,
            DIN => \N__3467\,
            DOUT => \N__3466\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3468\,
            PADOUT => \N__3467\,
            PADIN => \N__3466\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2627\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3459\,
            DIN => \N__3458\,
            DOUT => \N__3457\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3459\,
            PADOUT => \N__3458\,
            PADIN => \N__3457\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2111\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3450\,
            DIN => \N__3449\,
            DOUT => \N__3448\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3450\,
            PADOUT => \N__3449\,
            PADIN => \N__3448\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2168\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3441\,
            DIN => \N__3440\,
            DOUT => \N__3439\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3441\,
            PADOUT => \N__3440\,
            PADIN => \N__3439\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2204\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3432\,
            DIN => \N__3431\,
            DOUT => \N__3430\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3432\,
            PADOUT => \N__3431\,
            PADIN => \N__3430\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2936\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3423\,
            DIN => \N__3422\,
            DOUT => \N__3421\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3423\,
            PADOUT => \N__3422\,
            PADIN => \N__3421\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2009\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3414\,
            DIN => \N__3413\,
            DOUT => \N__3412\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3414\,
            PADOUT => \N__3413\,
            PADIN => \N__3412\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1961\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3405\,
            DIN => \N__3404\,
            DOUT => \N__3403\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3405\,
            PADOUT => \N__3404\,
            PADIN => \N__3403\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1556\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3396\,
            DIN => \N__3395\,
            DOUT => \N__3394\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3396\,
            PADOUT => \N__3395\,
            PADIN => \N__3394\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \trigger_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3387\,
            DIN => \N__3386\,
            DOUT => \N__3385\,
            PACKAGEPIN => trigger_wire
        );

    \trigger_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3387\,
            PADOUT => \N__3386\,
            PADIN => \N__3385\,
            CLOCKENABLE => 'H',
            DIN0 => trigger_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \usb_tx_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3378\,
            DIN => \N__3377\,
            DOUT => \N__3376\,
            PACKAGEPIN => usb_tx_wire
        );

    \usb_tx_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3378\,
            PADOUT => \N__3377\,
            PADIN => \N__3376\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1406\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__775\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3356\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3356\,
            I => \N__3352\
        );

    \I__773\ : InMux
    port map (
            O => \N__3355\,
            I => \N__3348\
        );

    \I__772\ : Span4Mux_h
    port map (
            O => \N__3352\,
            I => \N__3345\
        );

    \I__771\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3342\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3348\,
            I => \btn_cond.M_ctr_qZ0Z_13\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__3345\,
            I => \btn_cond.M_ctr_qZ0Z_13\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3342\,
            I => \btn_cond.M_ctr_qZ0Z_13\
        );

    \I__767\ : InMux
    port map (
            O => \N__3335\,
            I => \btn_cond.un1_M_ctr_q_cry_12\
        );

    \I__766\ : InMux
    port map (
            O => \N__3332\,
            I => \N__3328\
        );

    \I__765\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3325\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3328\,
            I => \N__3322\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3325\,
            I => \N__3316\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__3322\,
            I => \N__3316\
        );

    \I__761\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3313\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__3316\,
            I => \btn_cond.M_ctr_qZ0Z_14\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3313\,
            I => \btn_cond.M_ctr_qZ0Z_14\
        );

    \I__758\ : InMux
    port map (
            O => \N__3308\,
            I => \btn_cond.un1_M_ctr_q_cry_13\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__3305\,
            I => \N__3301\
        );

    \I__756\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3297\
        );

    \I__755\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3294\
        );

    \I__754\ : InMux
    port map (
            O => \N__3300\,
            I => \N__3291\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3297\,
            I => \btn_cond.M_ctr_qZ0Z_15\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3294\,
            I => \btn_cond.M_ctr_qZ0Z_15\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3291\,
            I => \btn_cond.M_ctr_qZ0Z_15\
        );

    \I__750\ : InMux
    port map (
            O => \N__3284\,
            I => \btn_cond.un1_M_ctr_q_cry_14\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__3281\,
            I => \N__3277\
        );

    \I__748\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3271\
        );

    \I__747\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3271\
        );

    \I__746\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3268\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3271\,
            I => \N__3265\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3268\,
            I => \btn_cond.M_ctr_qZ0Z_16\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__3265\,
            I => \btn_cond.M_ctr_qZ0Z_16\
        );

    \I__742\ : InMux
    port map (
            O => \N__3260\,
            I => \bfn_18_29_0_\
        );

    \I__741\ : InMux
    port map (
            O => \N__3257\,
            I => \N__3250\
        );

    \I__740\ : InMux
    port map (
            O => \N__3256\,
            I => \N__3250\
        );

    \I__739\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3247\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3250\,
            I => \N__3244\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3247\,
            I => \btn_cond.M_ctr_qZ0Z_17\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__3244\,
            I => \btn_cond.M_ctr_qZ0Z_17\
        );

    \I__735\ : InMux
    port map (
            O => \N__3239\,
            I => \btn_cond.un1_M_ctr_q_cry_16\
        );

    \I__734\ : InMux
    port map (
            O => \N__3236\,
            I => \N__3231\
        );

    \I__733\ : InMux
    port map (
            O => \N__3235\,
            I => \N__3226\
        );

    \I__732\ : InMux
    port map (
            O => \N__3234\,
            I => \N__3226\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3231\,
            I => \btn_cond.M_ctr_qZ0Z_18\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3226\,
            I => \btn_cond.M_ctr_qZ0Z_18\
        );

    \I__729\ : InMux
    port map (
            O => \N__3221\,
            I => \btn_cond.un1_M_ctr_q_cry_17\
        );

    \I__728\ : InMux
    port map (
            O => \N__3218\,
            I => \btn_cond.un1_M_ctr_q_cry_18\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__3215\,
            I => \N__3211\
        );

    \I__726\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3207\
        );

    \I__725\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3202\
        );

    \I__724\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3202\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3207\,
            I => \btn_cond.M_ctr_qZ0Z_19\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3202\,
            I => \btn_cond.M_ctr_qZ0Z_19\
        );

    \I__721\ : ClkMux
    port map (
            O => \N__3197\,
            I => \N__3149\
        );

    \I__720\ : ClkMux
    port map (
            O => \N__3196\,
            I => \N__3149\
        );

    \I__719\ : ClkMux
    port map (
            O => \N__3195\,
            I => \N__3149\
        );

    \I__718\ : ClkMux
    port map (
            O => \N__3194\,
            I => \N__3149\
        );

    \I__717\ : ClkMux
    port map (
            O => \N__3193\,
            I => \N__3149\
        );

    \I__716\ : ClkMux
    port map (
            O => \N__3192\,
            I => \N__3149\
        );

    \I__715\ : ClkMux
    port map (
            O => \N__3191\,
            I => \N__3149\
        );

    \I__714\ : ClkMux
    port map (
            O => \N__3190\,
            I => \N__3149\
        );

    \I__713\ : ClkMux
    port map (
            O => \N__3189\,
            I => \N__3149\
        );

    \I__712\ : ClkMux
    port map (
            O => \N__3188\,
            I => \N__3149\
        );

    \I__711\ : ClkMux
    port map (
            O => \N__3187\,
            I => \N__3149\
        );

    \I__710\ : ClkMux
    port map (
            O => \N__3186\,
            I => \N__3149\
        );

    \I__709\ : ClkMux
    port map (
            O => \N__3185\,
            I => \N__3149\
        );

    \I__708\ : ClkMux
    port map (
            O => \N__3184\,
            I => \N__3149\
        );

    \I__707\ : ClkMux
    port map (
            O => \N__3183\,
            I => \N__3149\
        );

    \I__706\ : ClkMux
    port map (
            O => \N__3182\,
            I => \N__3149\
        );

    \I__705\ : GlobalMux
    port map (
            O => \N__3149\,
            I => \N__3146\
        );

    \I__704\ : gio2CtrlBuf
    port map (
            O => \N__3146\,
            I => clk_c_g
        );

    \I__703\ : SRMux
    port map (
            O => \N__3143\,
            I => \N__3134\
        );

    \I__702\ : SRMux
    port map (
            O => \N__3142\,
            I => \N__3134\
        );

    \I__701\ : SRMux
    port map (
            O => \N__3141\,
            I => \N__3134\
        );

    \I__700\ : GlobalMux
    port map (
            O => \N__3134\,
            I => \N__3131\
        );

    \I__699\ : gio2CtrlBuf
    port map (
            O => \N__3131\,
            I => \btn_cond.M_sync_out_i_g_0\
        );

    \I__698\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3123\
        );

    \I__697\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3120\
        );

    \I__696\ : InMux
    port map (
            O => \N__3126\,
            I => \N__3117\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3123\,
            I => \btn_cond.M_ctr_qZ0Z_5\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3120\,
            I => \btn_cond.M_ctr_qZ0Z_5\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3117\,
            I => \btn_cond.M_ctr_qZ0Z_5\
        );

    \I__692\ : InMux
    port map (
            O => \N__3110\,
            I => \btn_cond.un1_M_ctr_q_cry_4\
        );

    \I__691\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3102\
        );

    \I__690\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3099\
        );

    \I__689\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3096\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3102\,
            I => \btn_cond.M_ctr_qZ0Z_6\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3099\,
            I => \btn_cond.M_ctr_qZ0Z_6\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3096\,
            I => \btn_cond.M_ctr_qZ0Z_6\
        );

    \I__685\ : InMux
    port map (
            O => \N__3089\,
            I => \btn_cond.un1_M_ctr_q_cry_5\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__3086\,
            I => \N__3081\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__3085\,
            I => \N__3078\
        );

    \I__682\ : InMux
    port map (
            O => \N__3084\,
            I => \N__3075\
        );

    \I__681\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3072\
        );

    \I__680\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3069\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3075\,
            I => \N__3064\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3072\,
            I => \N__3064\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3069\,
            I => \btn_cond.M_ctr_qZ0Z_7\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__3064\,
            I => \btn_cond.M_ctr_qZ0Z_7\
        );

    \I__675\ : InMux
    port map (
            O => \N__3059\,
            I => \btn_cond.un1_M_ctr_q_cry_6\
        );

    \I__674\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3052\
        );

    \I__673\ : InMux
    port map (
            O => \N__3055\,
            I => \N__3048\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3052\,
            I => \N__3045\
        );

    \I__671\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3042\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3048\,
            I => \btn_cond.M_ctr_qZ0Z_8\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__3045\,
            I => \btn_cond.M_ctr_qZ0Z_8\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3042\,
            I => \btn_cond.M_ctr_qZ0Z_8\
        );

    \I__667\ : InMux
    port map (
            O => \N__3035\,
            I => \bfn_18_28_0_\
        );

    \I__666\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3027\
        );

    \I__665\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3024\
        );

    \I__664\ : InMux
    port map (
            O => \N__3030\,
            I => \N__3021\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3027\,
            I => \btn_cond.M_ctr_qZ0Z_9\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3024\,
            I => \btn_cond.M_ctr_qZ0Z_9\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3021\,
            I => \btn_cond.M_ctr_qZ0Z_9\
        );

    \I__660\ : InMux
    port map (
            O => \N__3014\,
            I => \btn_cond.un1_M_ctr_q_cry_8\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__3011\,
            I => \N__3007\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__3010\,
            I => \N__3003\
        );

    \I__657\ : InMux
    port map (
            O => \N__3007\,
            I => \N__3000\
        );

    \I__656\ : InMux
    port map (
            O => \N__3006\,
            I => \N__2997\
        );

    \I__655\ : InMux
    port map (
            O => \N__3003\,
            I => \N__2994\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3000\,
            I => \N__2991\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__2997\,
            I => \btn_cond.M_ctr_qZ0Z_10\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__2994\,
            I => \btn_cond.M_ctr_qZ0Z_10\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__2991\,
            I => \btn_cond.M_ctr_qZ0Z_10\
        );

    \I__650\ : InMux
    port map (
            O => \N__2984\,
            I => \btn_cond.un1_M_ctr_q_cry_9\
        );

    \I__649\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2976\
        );

    \I__648\ : InMux
    port map (
            O => \N__2980\,
            I => \N__2973\
        );

    \I__647\ : InMux
    port map (
            O => \N__2979\,
            I => \N__2970\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__2976\,
            I => \btn_cond.M_ctr_qZ0Z_11\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__2973\,
            I => \btn_cond.M_ctr_qZ0Z_11\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__2970\,
            I => \btn_cond.M_ctr_qZ0Z_11\
        );

    \I__643\ : InMux
    port map (
            O => \N__2963\,
            I => \btn_cond.un1_M_ctr_q_cry_10\
        );

    \I__642\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2955\
        );

    \I__641\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2952\
        );

    \I__640\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2949\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__2955\,
            I => \btn_cond.M_ctr_qZ0Z_12\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__2952\,
            I => \btn_cond.M_ctr_qZ0Z_12\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__2949\,
            I => \btn_cond.M_ctr_qZ0Z_12\
        );

    \I__636\ : InMux
    port map (
            O => \N__2942\,
            I => \btn_cond.un1_M_ctr_q_cry_11\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__2939\,
            I => \un1_M_count_q_ac0_5_m2_0_a2_3_cascade_\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__2936\,
            I => \N__2933\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__632\ : IoSpan4Mux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__631\ : Span4Mux_s2_h
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__2924\,
            I => \N__2920\
        );

    \I__629\ : InMux
    port map (
            O => \N__2923\,
            I => \N__2917\
        );

    \I__628\ : Span12Mux_v
    port map (
            O => \N__2920\,
            I => \N__2913\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__2917\,
            I => \N__2910\
        );

    \I__626\ : InMux
    port map (
            O => \N__2916\,
            I => \N__2907\
        );

    \I__625\ : Span12Mux_h
    port map (
            O => \N__2913\,
            I => \N__2903\
        );

    \I__624\ : Span4Mux_h
    port map (
            O => \N__2910\,
            I => \N__2900\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__2907\,
            I => \N__2897\
        );

    \I__622\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2894\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__2903\,
            I => led_c_4
        );

    \I__620\ : Odrv4
    port map (
            O => \N__2900\,
            I => led_c_4
        );

    \I__619\ : Odrv4
    port map (
            O => \N__2897\,
            I => led_c_4
        );

    \I__618\ : LocalMux
    port map (
            O => \N__2894\,
            I => led_c_4
        );

    \I__617\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2879\
        );

    \I__616\ : InMux
    port map (
            O => \N__2884\,
            I => \N__2876\
        );

    \I__615\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2873\
        );

    \I__614\ : InMux
    port map (
            O => \N__2882\,
            I => \N__2870\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__2879\,
            I => \N__2865\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2876\,
            I => \N__2865\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__2873\,
            I => btn_cond_out_16_5
        );

    \I__610\ : LocalMux
    port map (
            O => \N__2870\,
            I => btn_cond_out_16_5
        );

    \I__609\ : Odrv4
    port map (
            O => \N__2865\,
            I => btn_cond_out_16_5
        );

    \I__608\ : InMux
    port map (
            O => \N__2858\,
            I => \N__2855\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__2855\,
            I => \N__2848\
        );

    \I__606\ : InMux
    port map (
            O => \N__2854\,
            I => \N__2843\
        );

    \I__605\ : InMux
    port map (
            O => \N__2853\,
            I => \N__2843\
        );

    \I__604\ : InMux
    port map (
            O => \N__2852\,
            I => \N__2840\
        );

    \I__603\ : InMux
    port map (
            O => \N__2851\,
            I => \N__2837\
        );

    \I__602\ : Span4Mux_h
    port map (
            O => \N__2848\,
            I => \N__2832\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__2843\,
            I => \N__2832\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__2840\,
            I => \N__2827\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__2837\,
            I => \N__2827\
        );

    \I__598\ : Odrv4
    port map (
            O => \N__2832\,
            I => btn_cond_out_16_4
        );

    \I__597\ : Odrv12
    port map (
            O => \N__2827\,
            I => btn_cond_out_16_4
        );

    \I__596\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2816\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__2821\,
            I => \N__2813\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__2820\,
            I => \N__2808\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__2819\,
            I => \N__2805\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__2816\,
            I => \N__2802\
        );

    \I__591\ : InMux
    port map (
            O => \N__2813\,
            I => \N__2799\
        );

    \I__590\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2796\
        );

    \I__589\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2789\
        );

    \I__588\ : InMux
    port map (
            O => \N__2808\,
            I => \N__2789\
        );

    \I__587\ : InMux
    port map (
            O => \N__2805\,
            I => \N__2789\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__2802\,
            I => \click_dtct_M_last_q\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__2799\,
            I => \click_dtct_M_last_q\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__2796\,
            I => \click_dtct_M_last_q\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__2789\,
            I => \click_dtct_M_last_q\
        );

    \I__582\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2776\
        );

    \I__581\ : InMux
    port map (
            O => \N__2779\,
            I => \N__2770\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__2776\,
            I => \N__2767\
        );

    \I__579\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2762\
        );

    \I__578\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2762\
        );

    \I__577\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2759\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__2770\,
            I => btn_cond_out_17
        );

    \I__575\ : Odrv4
    port map (
            O => \N__2767\,
            I => btn_cond_out_17
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2762\,
            I => btn_cond_out_17
        );

    \I__573\ : LocalMux
    port map (
            O => \N__2759\,
            I => btn_cond_out_17
        );

    \I__572\ : InMux
    port map (
            O => \N__2750\,
            I => \N__2745\
        );

    \I__571\ : InMux
    port map (
            O => \N__2749\,
            I => \N__2740\
        );

    \I__570\ : InMux
    port map (
            O => \N__2748\,
            I => \N__2740\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__2745\,
            I => click_dtct_out8
        );

    \I__568\ : LocalMux
    port map (
            O => \N__2740\,
            I => click_dtct_out8
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__2735\,
            I => \N__2729\
        );

    \I__566\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2721\
        );

    \I__565\ : InMux
    port map (
            O => \N__2733\,
            I => \N__2721\
        );

    \I__564\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2721\
        );

    \I__563\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2716\
        );

    \I__562\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2716\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__2721\,
            I => click_dtct_out3
        );

    \I__560\ : LocalMux
    port map (
            O => \N__2716\,
            I => click_dtct_out3
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__2711\,
            I => \click_dtct_out8_cascade_\
        );

    \I__558\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2699\
        );

    \I__557\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2694\
        );

    \I__556\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2694\
        );

    \I__555\ : InMux
    port map (
            O => \N__2705\,
            I => \N__2687\
        );

    \I__554\ : InMux
    port map (
            O => \N__2704\,
            I => \N__2687\
        );

    \I__553\ : InMux
    port map (
            O => \N__2703\,
            I => \N__2687\
        );

    \I__552\ : SRMux
    port map (
            O => \N__2702\,
            I => \N__2684\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__2699\,
            I => \N__2675\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__2694\,
            I => \N__2675\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2687\,
            I => \N__2670\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2684\,
            I => \N__2670\
        );

    \I__547\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2663\
        );

    \I__546\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2656\
        );

    \I__545\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2656\
        );

    \I__544\ : InMux
    port map (
            O => \N__2680\,
            I => \N__2656\
        );

    \I__543\ : Span4Mux_v
    port map (
            O => \N__2675\,
            I => \N__2651\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__2670\,
            I => \N__2651\
        );

    \I__541\ : InMux
    port map (
            O => \N__2669\,
            I => \N__2648\
        );

    \I__540\ : InMux
    port map (
            O => \N__2668\,
            I => \N__2645\
        );

    \I__539\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2640\
        );

    \I__538\ : InMux
    port map (
            O => \N__2666\,
            I => \N__2640\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__2663\,
            I => \uart_tx_N_186_1\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2656\,
            I => \uart_tx_N_186_1\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__2651\,
            I => \uart_tx_N_186_1\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__2648\,
            I => \uart_tx_N_186_1\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2645\,
            I => \uart_tx_N_186_1\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2640\,
            I => \uart_tx_N_186_1\
        );

    \I__531\ : IoInMux
    port map (
            O => \N__2627\,
            I => \N__2624\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__2624\,
            I => \N__2621\
        );

    \I__529\ : IoSpan4Mux
    port map (
            O => \N__2621\,
            I => \N__2618\
        );

    \I__528\ : Span4Mux_s3_h
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__527\ : Sp12to4
    port map (
            O => \N__2615\,
            I => \N__2611\
        );

    \I__526\ : InMux
    port map (
            O => \N__2614\,
            I => \N__2608\
        );

    \I__525\ : Span12Mux_h
    port map (
            O => \N__2611\,
            I => \N__2605\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__2608\,
            I => \N__2602\
        );

    \I__523\ : Span12Mux_v
    port map (
            O => \N__2605\,
            I => \N__2596\
        );

    \I__522\ : Span4Mux_h
    port map (
            O => \N__2602\,
            I => \N__2593\
        );

    \I__521\ : InMux
    port map (
            O => \N__2601\,
            I => \N__2590\
        );

    \I__520\ : InMux
    port map (
            O => \N__2600\,
            I => \N__2587\
        );

    \I__519\ : InMux
    port map (
            O => \N__2599\,
            I => \N__2584\
        );

    \I__518\ : Odrv12
    port map (
            O => \N__2596\,
            I => led_c_0
        );

    \I__517\ : Odrv4
    port map (
            O => \N__2593\,
            I => led_c_0
        );

    \I__516\ : LocalMux
    port map (
            O => \N__2590\,
            I => led_c_0
        );

    \I__515\ : LocalMux
    port map (
            O => \N__2587\,
            I => led_c_0
        );

    \I__514\ : LocalMux
    port map (
            O => \N__2584\,
            I => led_c_0
        );

    \I__513\ : SRMux
    port map (
            O => \N__2573\,
            I => \N__2568\
        );

    \I__512\ : SRMux
    port map (
            O => \N__2572\,
            I => \N__2565\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__2571\,
            I => \N__2560\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__2568\,
            I => \N__2557\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__2565\,
            I => \N__2554\
        );

    \I__508\ : SRMux
    port map (
            O => \N__2564\,
            I => \N__2551\
        );

    \I__507\ : InMux
    port map (
            O => \N__2563\,
            I => \N__2548\
        );

    \I__506\ : InMux
    port map (
            O => \N__2560\,
            I => \N__2545\
        );

    \I__505\ : Span4Mux_v
    port map (
            O => \N__2557\,
            I => \N__2542\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__2554\,
            I => \N__2539\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2551\,
            I => \N__2536\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__2548\,
            I => \N__2533\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2545\,
            I => \N__2530\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__2542\,
            I => \M_reset_cond_out_0\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__2539\,
            I => \M_reset_cond_out_0\
        );

    \I__498\ : Odrv12
    port map (
            O => \N__2536\,
            I => \M_reset_cond_out_0\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__2533\,
            I => \M_reset_cond_out_0\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__2530\,
            I => \M_reset_cond_out_0\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__2519\,
            I => \N__2515\
        );

    \I__494\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2512\
        );

    \I__493\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2509\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2512\,
            I => \btn_cond.M_btn_cond_out_i_0\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2509\,
            I => \btn_cond.M_btn_cond_out_i_0\
        );

    \I__490\ : InMux
    port map (
            O => \N__2504\,
            I => \N__2499\
        );

    \I__489\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2496\
        );

    \I__488\ : InMux
    port map (
            O => \N__2502\,
            I => \N__2493\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__2499\,
            I => \btn_cond.M_ctr_qZ0Z_0\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2496\,
            I => \btn_cond.M_ctr_qZ0Z_0\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__2493\,
            I => \btn_cond.M_ctr_qZ0Z_0\
        );

    \I__484\ : InMux
    port map (
            O => \N__2486\,
            I => \N__2481\
        );

    \I__483\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2478\
        );

    \I__482\ : InMux
    port map (
            O => \N__2484\,
            I => \N__2475\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2481\,
            I => \btn_cond.M_ctr_qZ0Z_1\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2478\,
            I => \btn_cond.M_ctr_qZ0Z_1\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2475\,
            I => \btn_cond.M_ctr_qZ0Z_1\
        );

    \I__478\ : InMux
    port map (
            O => \N__2468\,
            I => \btn_cond.un1_M_ctr_q_cry_0\
        );

    \I__477\ : InMux
    port map (
            O => \N__2465\,
            I => \N__2460\
        );

    \I__476\ : InMux
    port map (
            O => \N__2464\,
            I => \N__2457\
        );

    \I__475\ : InMux
    port map (
            O => \N__2463\,
            I => \N__2454\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2460\,
            I => \N__2451\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__2457\,
            I => \btn_cond.M_ctr_qZ0Z_2\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2454\,
            I => \btn_cond.M_ctr_qZ0Z_2\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__2451\,
            I => \btn_cond.M_ctr_qZ0Z_2\
        );

    \I__470\ : InMux
    port map (
            O => \N__2444\,
            I => \btn_cond.un1_M_ctr_q_cry_1\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__2441\,
            I => \N__2437\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__2440\,
            I => \N__2433\
        );

    \I__467\ : InMux
    port map (
            O => \N__2437\,
            I => \N__2430\
        );

    \I__466\ : InMux
    port map (
            O => \N__2436\,
            I => \N__2427\
        );

    \I__465\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2424\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2430\,
            I => \N__2421\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2427\,
            I => \btn_cond.M_ctr_qZ0Z_3\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2424\,
            I => \btn_cond.M_ctr_qZ0Z_3\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__2421\,
            I => \btn_cond.M_ctr_qZ0Z_3\
        );

    \I__460\ : InMux
    port map (
            O => \N__2414\,
            I => \btn_cond.un1_M_ctr_q_cry_2\
        );

    \I__459\ : InMux
    port map (
            O => \N__2411\,
            I => \N__2406\
        );

    \I__458\ : InMux
    port map (
            O => \N__2410\,
            I => \N__2403\
        );

    \I__457\ : InMux
    port map (
            O => \N__2409\,
            I => \N__2400\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2406\,
            I => \btn_cond.M_ctr_qZ0Z_4\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2403\,
            I => \btn_cond.M_ctr_qZ0Z_4\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2400\,
            I => \btn_cond.M_ctr_qZ0Z_4\
        );

    \I__453\ : InMux
    port map (
            O => \N__2393\,
            I => \btn_cond.un1_M_ctr_q_cry_3\
        );

    \I__452\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2387\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2387\,
            I => \reset_cond.M_stage_qZ0Z_2\
        );

    \I__450\ : InMux
    port map (
            O => \N__2384\,
            I => \N__2372\
        );

    \I__449\ : InMux
    port map (
            O => \N__2383\,
            I => \N__2372\
        );

    \I__448\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2372\
        );

    \I__447\ : InMux
    port map (
            O => \N__2381\,
            I => \N__2372\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2372\,
            I => \N__2369\
        );

    \I__445\ : Span4Mux_v
    port map (
            O => \N__2369\,
            I => \N__2366\
        );

    \I__444\ : Sp12to4
    port map (
            O => \N__2366\,
            I => \N__2363\
        );

    \I__443\ : Span12Mux_h
    port map (
            O => \N__2363\,
            I => \N__2360\
        );

    \I__442\ : Span12Mux_v
    port map (
            O => \N__2360\,
            I => \N__2357\
        );

    \I__441\ : Odrv12
    port map (
            O => \N__2357\,
            I => rst_n_c
        );

    \I__440\ : InMux
    port map (
            O => \N__2354\,
            I => \N__2351\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2351\,
            I => \reset_cond.M_stage_qZ0Z_0\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__437\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2341\
        );

    \I__436\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2338\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2341\,
            I => \N__2335\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2338\,
            I => \uart_tx.N_186_1_i\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__2335\,
            I => \uart_tx.N_186_1_i\
        );

    \I__432\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2327\,
            I => \click_dtct_M_count_d6_0_1\
        );

    \I__430\ : InMux
    port map (
            O => \N__2324\,
            I => \N__2321\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2321\,
            I => \N__2311\
        );

    \I__428\ : InMux
    port map (
            O => \N__2320\,
            I => \N__2306\
        );

    \I__427\ : InMux
    port map (
            O => \N__2319\,
            I => \N__2306\
        );

    \I__426\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2299\
        );

    \I__425\ : InMux
    port map (
            O => \N__2317\,
            I => \N__2299\
        );

    \I__424\ : InMux
    port map (
            O => \N__2316\,
            I => \N__2299\
        );

    \I__423\ : InMux
    port map (
            O => \N__2315\,
            I => \N__2296\
        );

    \I__422\ : InMux
    port map (
            O => \N__2314\,
            I => \N__2293\
        );

    \I__421\ : Odrv4
    port map (
            O => \N__2311\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__2306\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2299\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2296\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2293\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__416\ : InMux
    port map (
            O => \N__2282\,
            I => \N__2278\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__2281\,
            I => \N__2272\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2278\,
            I => \N__2269\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2277\,
            I => \N__2266\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__2276\,
            I => \N__2263\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__2275\,
            I => \N__2260\
        );

    \I__410\ : InMux
    port map (
            O => \N__2272\,
            I => \N__2253\
        );

    \I__409\ : Span4Mux_v
    port map (
            O => \N__2269\,
            I => \N__2250\
        );

    \I__408\ : InMux
    port map (
            O => \N__2266\,
            I => \N__2245\
        );

    \I__407\ : InMux
    port map (
            O => \N__2263\,
            I => \N__2245\
        );

    \I__406\ : InMux
    port map (
            O => \N__2260\,
            I => \N__2238\
        );

    \I__405\ : InMux
    port map (
            O => \N__2259\,
            I => \N__2238\
        );

    \I__404\ : InMux
    port map (
            O => \N__2258\,
            I => \N__2238\
        );

    \I__403\ : InMux
    port map (
            O => \N__2257\,
            I => \N__2235\
        );

    \I__402\ : InMux
    port map (
            O => \N__2256\,
            I => \N__2232\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2253\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__400\ : Odrv4
    port map (
            O => \N__2250\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2245\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2238\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2235\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2232\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__2219\,
            I => \uart_tx_N_186_1_cascade_\
        );

    \I__394\ : InMux
    port map (
            O => \N__2216\,
            I => \N__2212\
        );

    \I__393\ : InMux
    port map (
            O => \N__2215\,
            I => \N__2209\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2212\,
            I => \un1_M_count_q_ac0_out\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2209\,
            I => \un1_M_count_q_ac0_out\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__2204\,
            I => \N__2201\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2201\,
            I => \N__2198\
        );

    \I__388\ : Span12Mux_s3_h
    port map (
            O => \N__2198\,
            I => \N__2195\
        );

    \I__387\ : Span12Mux_h
    port map (
            O => \N__2195\,
            I => \N__2192\
        );

    \I__386\ : Span12Mux_v
    port map (
            O => \N__2192\,
            I => \N__2186\
        );

    \I__385\ : InMux
    port map (
            O => \N__2191\,
            I => \N__2183\
        );

    \I__384\ : InMux
    port map (
            O => \N__2190\,
            I => \N__2180\
        );

    \I__383\ : InMux
    port map (
            O => \N__2189\,
            I => \N__2177\
        );

    \I__382\ : Odrv12
    port map (
            O => \N__2186\,
            I => led_c_3
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2183\,
            I => led_c_3
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2180\,
            I => led_c_3
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2177\,
            I => led_c_3
        );

    \I__378\ : IoInMux
    port map (
            O => \N__2168\,
            I => \N__2165\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2165\,
            I => \N__2162\
        );

    \I__376\ : IoSpan4Mux
    port map (
            O => \N__2162\,
            I => \N__2159\
        );

    \I__375\ : Span4Mux_s3_h
    port map (
            O => \N__2159\,
            I => \N__2156\
        );

    \I__374\ : Span4Mux_h
    port map (
            O => \N__2156\,
            I => \N__2153\
        );

    \I__373\ : Sp12to4
    port map (
            O => \N__2153\,
            I => \N__2150\
        );

    \I__372\ : Span12Mux_h
    port map (
            O => \N__2150\,
            I => \N__2145\
        );

    \I__371\ : InMux
    port map (
            O => \N__2149\,
            I => \N__2140\
        );

    \I__370\ : InMux
    port map (
            O => \N__2148\,
            I => \N__2137\
        );

    \I__369\ : Span12Mux_v
    port map (
            O => \N__2145\,
            I => \N__2134\
        );

    \I__368\ : InMux
    port map (
            O => \N__2144\,
            I => \N__2131\
        );

    \I__367\ : InMux
    port map (
            O => \N__2143\,
            I => \N__2128\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2140\,
            I => \N__2123\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2137\,
            I => \N__2123\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__2134\,
            I => led_c_2
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2131\,
            I => led_c_2
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2128\,
            I => led_c_2
        );

    \I__361\ : Odrv4
    port map (
            O => \N__2123\,
            I => led_c_2
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__2114\,
            I => \un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__2111\,
            I => \N__2108\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2108\,
            I => \N__2105\
        );

    \I__357\ : IoSpan4Mux
    port map (
            O => \N__2105\,
            I => \N__2102\
        );

    \I__356\ : Span4Mux_s3_h
    port map (
            O => \N__2102\,
            I => \N__2099\
        );

    \I__355\ : Sp12to4
    port map (
            O => \N__2099\,
            I => \N__2095\
        );

    \I__354\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2092\
        );

    \I__353\ : Span12Mux_h
    port map (
            O => \N__2095\,
            I => \N__2088\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2092\,
            I => \N__2085\
        );

    \I__351\ : CascadeMux
    port map (
            O => \N__2091\,
            I => \N__2081\
        );

    \I__350\ : Span12Mux_v
    port map (
            O => \N__2088\,
            I => \N__2077\
        );

    \I__349\ : Span4Mux_v
    port map (
            O => \N__2085\,
            I => \N__2074\
        );

    \I__348\ : InMux
    port map (
            O => \N__2084\,
            I => \N__2071\
        );

    \I__347\ : InMux
    port map (
            O => \N__2081\,
            I => \N__2066\
        );

    \I__346\ : InMux
    port map (
            O => \N__2080\,
            I => \N__2066\
        );

    \I__345\ : Odrv12
    port map (
            O => \N__2077\,
            I => led_c_1
        );

    \I__344\ : Odrv4
    port map (
            O => \N__2074\,
            I => led_c_1
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2071\,
            I => led_c_1
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2066\,
            I => led_c_1
        );

    \I__341\ : InMux
    port map (
            O => \N__2057\,
            I => \N__2054\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2054\,
            I => \N__2051\
        );

    \I__339\ : Odrv4
    port map (
            O => \N__2051\,
            I => \un1_M_count_q_ac0_5_m2_0_a2_3\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__2048\,
            I => \btn_cond.g0_13_cascade_\
        );

    \I__337\ : InMux
    port map (
            O => \N__2045\,
            I => \N__2042\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2042\,
            I => \btn_cond.g0_5\
        );

    \I__335\ : InMux
    port map (
            O => \N__2039\,
            I => \N__2036\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2036\,
            I => \btn_cond.g0_14\
        );

    \I__333\ : InMux
    port map (
            O => \N__2033\,
            I => \N__2030\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2030\,
            I => \btn_cond.g0_11\
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__2027\,
            I => \btn_cond.g0_16_cascade_\
        );

    \I__330\ : InMux
    port map (
            O => \N__2024\,
            I => \N__2021\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2021\,
            I => \btn_cond.g0_10\
        );

    \I__328\ : InMux
    port map (
            O => \N__2018\,
            I => \N__2015\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2015\,
            I => \reset_cond.M_stage_qZ0Z_1\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2012\,
            I => \un1_M_count_q_ac0_7_cascade_\
        );

    \I__325\ : IoInMux
    port map (
            O => \N__2009\,
            I => \N__2006\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2006\,
            I => \N__2003\
        );

    \I__323\ : IoSpan4Mux
    port map (
            O => \N__2003\,
            I => \N__2000\
        );

    \I__322\ : Sp12to4
    port map (
            O => \N__2000\,
            I => \N__1997\
        );

    \I__321\ : Span12Mux_s9_h
    port map (
            O => \N__1997\,
            I => \N__1994\
        );

    \I__320\ : Span12Mux_v
    port map (
            O => \N__1994\,
            I => \N__1991\
        );

    \I__319\ : Span12Mux_v
    port map (
            O => \N__1991\,
            I => \N__1984\
        );

    \I__318\ : InMux
    port map (
            O => \N__1990\,
            I => \N__1981\
        );

    \I__317\ : InMux
    port map (
            O => \N__1989\,
            I => \N__1978\
        );

    \I__316\ : InMux
    port map (
            O => \N__1988\,
            I => \N__1975\
        );

    \I__315\ : InMux
    port map (
            O => \N__1987\,
            I => \N__1972\
        );

    \I__314\ : Odrv12
    port map (
            O => \N__1984\,
            I => led_c_5
        );

    \I__313\ : LocalMux
    port map (
            O => \N__1981\,
            I => led_c_5
        );

    \I__312\ : LocalMux
    port map (
            O => \N__1978\,
            I => led_c_5
        );

    \I__311\ : LocalMux
    port map (
            O => \N__1975\,
            I => led_c_5
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1972\,
            I => led_c_5
        );

    \I__309\ : IoInMux
    port map (
            O => \N__1961\,
            I => \N__1958\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__1958\,
            I => \N__1955\
        );

    \I__307\ : Span12Mux_s6_h
    port map (
            O => \N__1955\,
            I => \N__1952\
        );

    \I__306\ : Span12Mux_v
    port map (
            O => \N__1952\,
            I => \N__1949\
        );

    \I__305\ : Span12Mux_v
    port map (
            O => \N__1949\,
            I => \N__1943\
        );

    \I__304\ : InMux
    port map (
            O => \N__1948\,
            I => \N__1940\
        );

    \I__303\ : InMux
    port map (
            O => \N__1947\,
            I => \N__1937\
        );

    \I__302\ : InMux
    port map (
            O => \N__1946\,
            I => \N__1934\
        );

    \I__301\ : Odrv12
    port map (
            O => \N__1943\,
            I => led_c_6
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1940\,
            I => led_c_6
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1937\,
            I => led_c_6
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1934\,
            I => led_c_6
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__1925\,
            I => \btn_cond_out_16_5_cascade_\
        );

    \I__296\ : InMux
    port map (
            O => \N__1922\,
            I => \N__1913\
        );

    \I__295\ : InMux
    port map (
            O => \N__1921\,
            I => \N__1913\
        );

    \I__294\ : InMux
    port map (
            O => \N__1920\,
            I => \N__1908\
        );

    \I__293\ : InMux
    port map (
            O => \N__1919\,
            I => \N__1908\
        );

    \I__292\ : InMux
    port map (
            O => \N__1918\,
            I => \N__1905\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1913\,
            I => click_dtct_out_d
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1908\,
            I => click_dtct_out_d
        );

    \I__289\ : LocalMux
    port map (
            O => \N__1905\,
            I => click_dtct_out_d
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__1898\,
            I => \btn_cond.out_17_8_cascade_\
        );

    \I__287\ : InMux
    port map (
            O => \N__1895\,
            I => \N__1892\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1892\,
            I => \btn_cond.out_17_6\
        );

    \I__285\ : InMux
    port map (
            O => \N__1889\,
            I => \N__1886\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1886\,
            I => \btn_cond.out_17_7\
        );

    \I__283\ : InMux
    port map (
            O => \N__1883\,
            I => \N__1875\
        );

    \I__282\ : InMux
    port map (
            O => \N__1882\,
            I => \N__1875\
        );

    \I__281\ : InMux
    port map (
            O => \N__1881\,
            I => \N__1872\
        );

    \I__280\ : InMux
    port map (
            O => \N__1880\,
            I => \N__1869\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1875\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1872\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__1869\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__276\ : InMux
    port map (
            O => \N__1862\,
            I => \N__1854\
        );

    \I__275\ : InMux
    port map (
            O => \N__1861\,
            I => \N__1851\
        );

    \I__274\ : InMux
    port map (
            O => \N__1860\,
            I => \N__1842\
        );

    \I__273\ : InMux
    port map (
            O => \N__1859\,
            I => \N__1842\
        );

    \I__272\ : InMux
    port map (
            O => \N__1858\,
            I => \N__1842\
        );

    \I__271\ : InMux
    port map (
            O => \N__1857\,
            I => \N__1842\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__1854\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1851\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1842\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__267\ : CascadeMux
    port map (
            O => \N__1835\,
            I => \uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_\
        );

    \I__266\ : InMux
    port map (
            O => \N__1832\,
            I => \N__1826\
        );

    \I__265\ : InMux
    port map (
            O => \N__1831\,
            I => \N__1820\
        );

    \I__264\ : InMux
    port map (
            O => \N__1830\,
            I => \N__1815\
        );

    \I__263\ : InMux
    port map (
            O => \N__1829\,
            I => \N__1815\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1826\,
            I => \N__1812\
        );

    \I__261\ : InMux
    port map (
            O => \N__1825\,
            I => \N__1805\
        );

    \I__260\ : InMux
    port map (
            O => \N__1824\,
            I => \N__1805\
        );

    \I__259\ : InMux
    port map (
            O => \N__1823\,
            I => \N__1805\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__1820\,
            I => \uart_tx.N_182_0\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1815\,
            I => \uart_tx.N_182_0\
        );

    \I__256\ : Odrv4
    port map (
            O => \N__1812\,
            I => \uart_tx.N_182_0\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1805\,
            I => \uart_tx.N_182_0\
        );

    \I__254\ : InMux
    port map (
            O => \N__1796\,
            I => \N__1789\
        );

    \I__253\ : InMux
    port map (
            O => \N__1795\,
            I => \N__1784\
        );

    \I__252\ : InMux
    port map (
            O => \N__1794\,
            I => \N__1784\
        );

    \I__251\ : InMux
    port map (
            O => \N__1793\,
            I => \N__1779\
        );

    \I__250\ : InMux
    port map (
            O => \N__1792\,
            I => \N__1779\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1789\,
            I => \uart_tx.M_bitCtr_qZ1Z_0\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1784\,
            I => \uart_tx.M_bitCtr_qZ1Z_0\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1779\,
            I => \uart_tx.M_bitCtr_qZ1Z_0\
        );

    \I__246\ : InMux
    port map (
            O => \N__1772\,
            I => \N__1769\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1769\,
            I => \uart_tx_N_185\
        );

    \I__244\ : CascadeMux
    port map (
            O => \N__1766\,
            I => \click_dtct_out3_cascade_\
        );

    \I__243\ : InMux
    port map (
            O => \N__1763\,
            I => \N__1760\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1760\,
            I => \uart_tx_N_187\
        );

    \I__241\ : InMux
    port map (
            O => \N__1757\,
            I => \N__1754\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__1754\,
            I => \un1_M_count_q_ac0_1\
        );

    \I__239\ : CascadeMux
    port map (
            O => \N__1751\,
            I => \un1_M_count_q_ac0_1_cascade_\
        );

    \I__238\ : CascadeMux
    port map (
            O => \N__1748\,
            I => \N__1745\
        );

    \I__237\ : InMux
    port map (
            O => \N__1745\,
            I => \N__1739\
        );

    \I__236\ : InMux
    port map (
            O => \N__1744\,
            I => \N__1739\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1739\,
            I => \un1_M_count_q_ac0_7\
        );

    \I__234\ : InMux
    port map (
            O => \N__1736\,
            I => \N__1732\
        );

    \I__233\ : InMux
    port map (
            O => \N__1735\,
            I => \N__1729\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1732\,
            I => \N__1726\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1729\,
            I => \uart_tx.M_ctr_qZ0Z_6\
        );

    \I__230\ : Odrv4
    port map (
            O => \N__1726\,
            I => \uart_tx.M_ctr_qZ0Z_6\
        );

    \I__229\ : InMux
    port map (
            O => \N__1721\,
            I => \N__1717\
        );

    \I__228\ : InMux
    port map (
            O => \N__1720\,
            I => \N__1714\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__1717\,
            I => \uart_tx.M_ctr_qZ1Z_4\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1714\,
            I => \uart_tx.M_ctr_qZ1Z_4\
        );

    \I__225\ : CascadeMux
    port map (
            O => \N__1709\,
            I => \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\
        );

    \I__224\ : InMux
    port map (
            O => \N__1706\,
            I => \N__1702\
        );

    \I__223\ : InMux
    port map (
            O => \N__1705\,
            I => \N__1699\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1702\,
            I => \uart_tx.M_ctr_qZ0Z_3\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1699\,
            I => \uart_tx.M_ctr_qZ0Z_3\
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__1694\,
            I => \uart_tx.N_182_0_cascade_\
        );

    \I__219\ : InMux
    port map (
            O => \N__1691\,
            I => \N__1688\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1688\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_2\
        );

    \I__217\ : InMux
    port map (
            O => \N__1685\,
            I => \N__1681\
        );

    \I__216\ : InMux
    port map (
            O => \N__1684\,
            I => \N__1678\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1681\,
            I => \N__1675\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1678\,
            I => \uart_tx.M_ctr_qZ0Z_2\
        );

    \I__213\ : Odrv4
    port map (
            O => \N__1675\,
            I => \uart_tx.M_ctr_qZ0Z_2\
        );

    \I__212\ : CascadeMux
    port map (
            O => \N__1670\,
            I => \N__1667\
        );

    \I__211\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1664\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1664\,
            I => \uart_tx.N_143_0\
        );

    \I__209\ : CascadeMux
    port map (
            O => \N__1661\,
            I => \uart_tx.N_143_0_cascade_\
        );

    \I__208\ : InMux
    port map (
            O => \N__1658\,
            I => \N__1654\
        );

    \I__207\ : InMux
    port map (
            O => \N__1657\,
            I => \N__1651\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1654\,
            I => \uart_tx.N_134_i\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__1651\,
            I => \uart_tx.N_134_i\
        );

    \I__204\ : CascadeMux
    port map (
            O => \N__1646\,
            I => \uart_tx.N_134_i_cascade_\
        );

    \I__203\ : InMux
    port map (
            O => \N__1643\,
            I => \N__1640\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1640\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_5\
        );

    \I__201\ : InMux
    port map (
            O => \N__1637\,
            I => \N__1633\
        );

    \I__200\ : InMux
    port map (
            O => \N__1636\,
            I => \N__1630\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1633\,
            I => \uart_tx.M_ctr_qZ1Z_5\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1630\,
            I => \uart_tx.M_ctr_qZ1Z_5\
        );

    \I__197\ : CascadeMux
    port map (
            O => \N__1625\,
            I => \M_btn_cond_out_0_cascade_\
        );

    \I__196\ : CEMux
    port map (
            O => \N__1622\,
            I => \N__1619\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1619\,
            I => \M_count_d6\
        );

    \I__194\ : InMux
    port map (
            O => \N__1616\,
            I => \uart_tx.un1_M_ctr_q_3_cry_0\
        );

    \I__193\ : InMux
    port map (
            O => \N__1613\,
            I => \uart_tx.un1_M_ctr_q_3_cry_1\
        );

    \I__192\ : InMux
    port map (
            O => \N__1610\,
            I => \uart_tx.un1_M_ctr_q_3_cry_2\
        );

    \I__191\ : InMux
    port map (
            O => \N__1607\,
            I => \uart_tx.un1_M_ctr_q_3_cry_3\
        );

    \I__190\ : InMux
    port map (
            O => \N__1604\,
            I => \uart_tx.un1_M_ctr_q_3_cry_4\
        );

    \I__189\ : InMux
    port map (
            O => \N__1601\,
            I => \uart_tx.un1_M_ctr_q_3_cry_5\
        );

    \I__188\ : CascadeMux
    port map (
            O => \N__1598\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__1595\,
            I => \N__1591\
        );

    \I__186\ : InMux
    port map (
            O => \N__1594\,
            I => \N__1588\
        );

    \I__185\ : InMux
    port map (
            O => \N__1591\,
            I => \N__1585\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1588\,
            I => \uart_tx.M_ctr_qZ0Z_0\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1585\,
            I => \uart_tx.M_ctr_qZ0Z_0\
        );

    \I__182\ : InMux
    port map (
            O => \N__1580\,
            I => \N__1576\
        );

    \I__181\ : InMux
    port map (
            O => \N__1579\,
            I => \N__1573\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1576\,
            I => \uart_tx.M_ctr_qZ1Z_1\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1573\,
            I => \uart_tx.M_ctr_qZ1Z_1\
        );

    \I__178\ : InMux
    port map (
            O => \N__1568\,
            I => \N__1565\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1565\,
            I => \uart_tx.M_savedData_qZ0Z_6\
        );

    \I__176\ : InMux
    port map (
            O => \N__1562\,
            I => \N__1559\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1559\,
            I => \uart_tx.M_savedData_qZ0Z_7\
        );

    \I__174\ : IoInMux
    port map (
            O => \N__1556\,
            I => \N__1553\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1553\,
            I => \N__1550\
        );

    \I__172\ : IoSpan4Mux
    port map (
            O => \N__1550\,
            I => \N__1547\
        );

    \I__171\ : Span4Mux_s0_v
    port map (
            O => \N__1547\,
            I => \N__1544\
        );

    \I__170\ : Sp12to4
    port map (
            O => \N__1544\,
            I => \N__1541\
        );

    \I__169\ : Span12Mux_s10_h
    port map (
            O => \N__1541\,
            I => \N__1538\
        );

    \I__168\ : Span12Mux_v
    port map (
            O => \N__1538\,
            I => \N__1535\
        );

    \I__167\ : Span12Mux_v
    port map (
            O => \N__1535\,
            I => \N__1530\
        );

    \I__166\ : InMux
    port map (
            O => \N__1534\,
            I => \N__1527\
        );

    \I__165\ : InMux
    port map (
            O => \N__1533\,
            I => \N__1524\
        );

    \I__164\ : Odrv12
    port map (
            O => \N__1530\,
            I => led_c_7
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1527\,
            I => led_c_7
        );

    \I__162\ : LocalMux
    port map (
            O => \N__1524\,
            I => led_c_7
        );

    \I__161\ : InMux
    port map (
            O => \N__1517\,
            I => \N__1514\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1514\,
            I => \un1_M_count_q_axbxc7_1\
        );

    \I__159\ : InMux
    port map (
            O => \N__1511\,
            I => \N__1508\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1508\,
            I => \N__1505\
        );

    \I__157\ : Span4Mux_v
    port map (
            O => \N__1505\,
            I => \N__1502\
        );

    \I__156\ : Sp12to4
    port map (
            O => \N__1502\,
            I => \N__1499\
        );

    \I__155\ : Span12Mux_h
    port map (
            O => \N__1499\,
            I => \N__1496\
        );

    \I__154\ : Span12Mux_v
    port map (
            O => \N__1496\,
            I => \N__1493\
        );

    \I__153\ : Odrv12
    port map (
            O => \N__1493\,
            I => trigger_c
        );

    \I__152\ : IoInMux
    port map (
            O => \N__1490\,
            I => \N__1487\
        );

    \I__151\ : LocalMux
    port map (
            O => \N__1487\,
            I => \btn_cond.sync.M_sync_out_i_0\
        );

    \I__150\ : InMux
    port map (
            O => \N__1484\,
            I => \N__1481\
        );

    \I__149\ : LocalMux
    port map (
            O => \N__1481\,
            I => \btn_cond.sync.M_pipe_qZ0Z_0\
        );

    \I__148\ : InMux
    port map (
            O => \N__1478\,
            I => \N__1475\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1475\,
            I => \btn_cond.sync.M_sync_out_0\
        );

    \I__146\ : CascadeMux
    port map (
            O => \N__1472\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_4_cascade_\
        );

    \I__145\ : InMux
    port map (
            O => \N__1469\,
            I => \N__1466\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__1466\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_5\
        );

    \I__143\ : InMux
    port map (
            O => \N__1463\,
            I => \N__1460\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__1460\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_2\
        );

    \I__141\ : CascadeMux
    port map (
            O => \N__1457\,
            I => \uart_tx.M_txReg_d_3_7_ns_1_cascade_\
        );

    \I__140\ : InMux
    port map (
            O => \N__1454\,
            I => \N__1451\
        );

    \I__139\ : LocalMux
    port map (
            O => \N__1451\,
            I => \uart_tx.M_txReg_q_RNOZ0Z_1\
        );

    \I__138\ : InMux
    port map (
            O => \N__1448\,
            I => \N__1445\
        );

    \I__137\ : LocalMux
    port map (
            O => \N__1445\,
            I => \uart_tx.M_txReg_d_3\
        );

    \I__136\ : InMux
    port map (
            O => \N__1442\,
            I => \N__1439\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__1439\,
            I => \uart_tx.M_savedData_qZ0Z_5\
        );

    \I__134\ : InMux
    port map (
            O => \N__1436\,
            I => \N__1433\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1433\,
            I => \uart_tx.M_savedData_qZ0Z_2\
        );

    \I__132\ : InMux
    port map (
            O => \N__1430\,
            I => \N__1427\
        );

    \I__131\ : LocalMux
    port map (
            O => \N__1427\,
            I => \uart_tx.M_savedData_qZ0Z_0\
        );

    \I__130\ : InMux
    port map (
            O => \N__1424\,
            I => \N__1421\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1421\,
            I => \uart_tx.M_savedData_qZ0Z_3\
        );

    \I__128\ : InMux
    port map (
            O => \N__1418\,
            I => \N__1415\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1415\,
            I => \uart_tx.M_savedData_qZ0Z_1\
        );

    \I__126\ : InMux
    port map (
            O => \N__1412\,
            I => \N__1409\
        );

    \I__125\ : LocalMux
    port map (
            O => \N__1409\,
            I => \uart_tx.M_savedData_qZ0Z_4\
        );

    \I__124\ : IoInMux
    port map (
            O => \N__1406\,
            I => \N__1403\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1403\,
            I => \N__1400\
        );

    \I__122\ : Span12Mux_s9_v
    port map (
            O => \N__1400\,
            I => \N__1397\
        );

    \I__121\ : Span12Mux_v
    port map (
            O => \N__1397\,
            I => \N__1394\
        );

    \I__120\ : Odrv12
    port map (
            O => \N__1394\,
            I => usb_tx_c
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_18_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_27_0_\
        );

    \IN_MUX_bfv_18_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \btn_cond.un1_M_ctr_q_cry_7\,
            carryinitout => \bfn_18_28_0_\
        );

    \IN_MUX_bfv_18_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \btn_cond.un1_M_ctr_q_cry_15\,
            carryinitout => \bfn_18_29_0_\
        );

    \btn_cond.sync.M_pipe_q_RNIJLM5_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1490\,
            GLOBALBUFFEROUTPUT => \btn_cond.M_sync_out_i_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111000110011"
        )
    port map (
            in0 => \N__1448\,
            in1 => \N__2282\,
            in2 => \_gnd_net_\,
            in3 => \N__2324\,
            lcout => usb_tx_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3182\,
            ce => 'H',
            sr => \N__2702\
        );

    \uart_tx.M_txReg_q_RNO_5_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__1568\,
            in1 => \N__1436\,
            in2 => \_gnd_net_\,
            in3 => \N__1857\,
            lcout => \uart_tx.M_txReg_q_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_2_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__1860\,
            in1 => \N__1562\,
            in2 => \_gnd_net_\,
            in3 => \N__1424\,
            lcout => \uart_tx.M_txReg_q_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_1_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__1442\,
            in1 => \N__1418\,
            in2 => \_gnd_net_\,
            in3 => \N__1859\,
            lcout => \uart_tx.M_txReg_q_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_4_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__1858\,
            in1 => \N__1412\,
            in2 => \_gnd_net_\,
            in3 => \N__1430\,
            lcout => OPEN,
            ltout => \uart_tx.M_txReg_q_RNOZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_3_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__1881\,
            in1 => \N__1794\,
            in2 => \N__1472\,
            in3 => \N__1469\,
            lcout => OPEN,
            ltout => \uart_tx.M_txReg_d_3_7_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_0_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__1795\,
            in1 => \N__1463\,
            in2 => \N__1457\,
            in3 => \N__1454\,
            lcout => \uart_tx.M_txReg_d_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_5_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1990\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_tx.M_savedData_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_2_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2144\,
            lcout => \uart_tx.M_savedData_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_0_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2614\,
            lcout => \uart_tx.M_savedData_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_3_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2191\,
            lcout => \uart_tx.M_savedData_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_1_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2098\,
            lcout => \uart_tx.M_savedData_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_4_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2923\,
            lcout => \uart_tx.M_savedData_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_6_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1948\,
            lcout => \uart_tx.M_savedData_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_7_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1534\,
            lcout => \uart_tx.M_savedData_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3184\,
            ce => \N__1622\,
            sr => \_gnd_net_\
        );

    \M_count_q_5_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__1922\,
            in1 => \N__1988\,
            in2 => \_gnd_net_\,
            in3 => \N__1744\,
            lcout => led_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3187\,
            ce => 'H',
            sr => \N__2573\
        );

    \M_count_q_7_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__1533\,
            in1 => \N__1946\,
            in2 => \N__1748\,
            in3 => \N__1517\,
            lcout => led_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3187\,
            ce => 'H',
            sr => \N__2573\
        );

    \M_count_q_2_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__2149\,
            in1 => \N__1921\,
            in2 => \_gnd_net_\,
            in3 => \N__1757\,
            lcout => led_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3187\,
            ce => 'H',
            sr => \N__2573\
        );

    \M_count_q_RNO_0_7_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1987\,
            in2 => \_gnd_net_\,
            in3 => \N__1918\,
            lcout => \un1_M_count_q_axbxc7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.sync.M_pipe_q_0_LC_16_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1511\,
            lcout => \btn_cond.sync.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.sync.M_pipe_q_RNIJLM5_1_LC_16_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1478\,
            lcout => \btn_cond.sync.M_sync_out_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.sync.M_pipe_q_1_LC_16_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1484\,
            lcout => \btn_cond.sync.M_sync_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_0_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2703\,
            in1 => \N__1594\,
            in2 => \N__2348\,
            in3 => \N__2344\,
            lcout => \uart_tx.M_ctr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_0\,
            clk => \N__3183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_1_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2706\,
            in1 => \N__1580\,
            in2 => \_gnd_net_\,
            in3 => \N__1616\,
            lcout => \uart_tx.M_ctr_qZ1Z_1\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_0\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_1\,
            clk => \N__3183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_2_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1684\,
            in2 => \_gnd_net_\,
            in3 => \N__1613\,
            lcout => \uart_tx.M_ctr_q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_1\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_3_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2707\,
            in1 => \N__1706\,
            in2 => \_gnd_net_\,
            in3 => \N__1610\,
            lcout => \uart_tx.M_ctr_qZ0Z_3\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_2\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_3\,
            clk => \N__3183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_4_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2704\,
            in1 => \N__1721\,
            in2 => \_gnd_net_\,
            in3 => \N__1607\,
            lcout => \uart_tx.M_ctr_qZ1Z_4\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_3\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_4\,
            clk => \N__3183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_5_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1637\,
            in2 => \_gnd_net_\,
            in3 => \N__1604\,
            lcout => \uart_tx.M_ctr_q_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_4\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_6_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1735\,
            in2 => \_gnd_net_\,
            in3 => \N__1601\,
            lcout => OPEN,
            ltout => \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_6_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__1658\,
            in1 => \N__2705\,
            in2 => \N__1598\,
            in3 => \N__1831\,
            lcout => \uart_tx.M_ctr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_2_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__1883\,
            in1 => \N__2682\,
            in2 => \N__1670\,
            in3 => \N__1862\,
            lcout => \uart_tx.M_bitCtr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNIGGUF1_0_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__1685\,
            in1 => \N__1636\,
            in2 => \N__1595\,
            in3 => \N__1579\,
            lcout => OPEN,
            ltout => \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNI3KTJ2_6_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__1736\,
            in1 => \N__1720\,
            in2 => \N__1709\,
            in3 => \N__1705\,
            lcout => \uart_tx.N_182_0\,
            ltout => \uart_tx.N_182_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_2_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__2680\,
            in1 => \N__1657\,
            in2 => \N__1694\,
            in3 => \N__1691\,
            lcout => \uart_tx.M_ctr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNIP5AF3_0_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2320\,
            in1 => \N__1796\,
            in2 => \N__2277\,
            in3 => \N__1829\,
            lcout => \uart_tx.N_143_0\,
            ltout => \uart_tx.N_143_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_1_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__2681\,
            in1 => \_gnd_net_\,
            in2 => \N__1661\,
            in3 => \N__1882\,
            lcout => \uart_tx.M_bitCtr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_0_1_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__2319\,
            in1 => \_gnd_net_\,
            in2 => \N__2276\,
            in3 => \_gnd_net_\,
            lcout => \uart_tx.N_134_i\,
            ltout => \uart_tx.N_134_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_5_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__1830\,
            in1 => \N__2708\,
            in2 => \N__1646\,
            in3 => \N__1643\,
            lcout => \uart_tx.M_ctr_qZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_1_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__1824\,
            in1 => \N__2318\,
            in2 => \N__2275\,
            in3 => \N__2563\,
            lcout => \uart_tx.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNICJ341_19_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2885\,
            in1 => \N__2852\,
            in2 => \_gnd_net_\,
            in3 => \N__2780\,
            lcout => OPEN,
            ltout => \M_btn_cond_out_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_RNIJC4S1_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2822\,
            in2 => \N__1625\,
            in3 => \N__2669\,
            lcout => \M_count_d6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNITA5V2_0_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2259\,
            in2 => \_gnd_net_\,
            in3 => \N__1823\,
            lcout => \uart_tx_N_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNITT1L_1_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__1880\,
            in1 => \N__1792\,
            in2 => \_gnd_net_\,
            in3 => \N__2258\,
            lcout => OPEN,
            ltout => \uart_tx.M_state_q_ns_0_a2_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNIUE4P3_2_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1861\,
            in1 => \N__1832\,
            in2 => \N__1835\,
            in3 => \N__2316\,
            lcout => \uart_tx_N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_0_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001011001000"
        )
    port map (
            in0 => \N__2317\,
            in1 => \N__1793\,
            in2 => \N__2281\,
            in3 => \N__1825\,
            lcout => \uart_tx.M_bitCtr_qZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_RNIUTK51_1_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2884\,
            in1 => \N__2851\,
            in2 => \N__2819\,
            in3 => \N__2773\,
            lcout => click_dtct_out3,
            ltout => \click_dtct_out3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_RNIE6EK8_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__2668\,
            in1 => \N__1772\,
            in2 => \N__1766\,
            in3 => \N__1763\,
            lcout => \click_dtct_M_count_d6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNI0H5P2_1_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__2084\,
            in1 => \N__2215\,
            in2 => \N__2820\,
            in3 => \N__2728\,
            lcout => \un1_M_count_q_ac0_1\,
            ltout => \un1_M_count_q_ac0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_3_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__2143\,
            in1 => \N__2190\,
            in2 => \N__1751\,
            in3 => \N__1919\,
            lcout => led_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3189\,
            ce => 'H',
            sr => \N__2572\
        );

    \M_count_q_RNIGFD24_4_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__2906\,
            in1 => \N__2811\,
            in2 => \N__2735\,
            in3 => \N__2057\,
            lcout => \un1_M_count_q_ac0_7\,
            ltout => \un1_M_count_q_ac0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_6_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__1920\,
            in1 => \N__1947\,
            in2 => \N__2012\,
            in3 => \N__1989\,
            lcout => led_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3189\,
            ce => 'H',
            sr => \N__2572\
        );

    \click_dtct.M_last_q_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2854\,
            in1 => \N__2883\,
            in2 => \_gnd_net_\,
            in3 => \N__2775\,
            lcout => \click_dtct_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIE6NB_0_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2463\,
            in1 => \N__2485\,
            in2 => \N__2440\,
            in3 => \N__2503\,
            lcout => btn_cond_out_16_5,
            ltout => \btn_cond_out_16_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click_dtct.M_last_q_RNIUTK51_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__2853\,
            in1 => \N__2812\,
            in2 => \N__1925\,
            in3 => \N__2774\,
            lcout => click_dtct_out_d,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIUMNB_4_LC_17_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3127\,
            in1 => \N__2410\,
            in2 => \N__3085\,
            in3 => \N__3106\,
            lcout => OPEN,
            ltout => \btn_cond.out_17_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIKBLL_10_LC_17_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1895\,
            in2 => \N__1898\,
            in3 => \N__1889\,
            lcout => btn_cond_out_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIQGM2_12_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3359\,
            in1 => \N__2959\,
            in2 => \N__3305\,
            in3 => \N__3332\,
            lcout => \btn_cond.out_17_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIS377_10_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3056\,
            in1 => \N__3031\,
            in2 => \N__3010\,
            in3 => \N__2980\,
            lcout => \btn_cond.out_17_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIE6NB_0_0_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__2465\,
            in1 => \N__2484\,
            in2 => \N__2441\,
            in3 => \N__2502\,
            lcout => \btn_cond.g0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIUMNB_0_4_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3105\,
            in1 => \N__3126\,
            in2 => \N__3086\,
            in3 => \N__2409\,
            lcout => \btn_cond.g0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIB6B1_12_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2958\,
            in2 => \_gnd_net_\,
            in3 => \N__3351\,
            lcout => \btn_cond.g0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIS377_0_10_LC_17_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3051\,
            in1 => \N__3030\,
            in2 => \N__3011\,
            in3 => \N__2979\,
            lcout => OPEN,
            ltout => \btn_cond.g0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIMKT9_14_LC_17_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__3300\,
            in1 => \N__3321\,
            in2 => \N__2048\,
            in3 => \N__2045\,
            lcout => OPEN,
            ltout => \btn_cond.g0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNICJ341_14_LC_17_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2039\,
            in1 => \N__2033\,
            in2 => \N__2027\,
            in3 => \N__2024\,
            lcout => \btn_cond.M_btn_cond_out_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIA1N2_0_19_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3256\,
            in1 => \N__3210\,
            in2 => \N__3281\,
            in3 => \N__3234\,
            lcout => \btn_cond.g0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \btn_cond.M_ctr_q_RNIA1N2_19_LC_17_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3235\,
            in1 => \N__3257\,
            in2 => \N__3215\,
            in3 => \N__3280\,
            lcout => btn_cond_out_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_2_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2383\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2018\,
            lcout => \reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_1_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2382\,
            in2 => \_gnd_net_\,
            in3 => \N__2354\,
            lcout => \reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_3_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2390\,
            lcout => \M_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_0_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2381\,
            lcout => \reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_1_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2257\,
            in2 => \_gnd_net_\,
            in3 => \N__2315\,
            lcout => \uart_tx.N_186_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_0_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001111"
        )
    port map (
            in0 => \N__2683\,
            in1 => \N__2750\,
            in2 => \N__2571\,
            in3 => \N__2330\,
            lcout => \uart_tx.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_1_1_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2314\,
            in2 => \_gnd_net_\,
            in3 => \N__2256\,
            lcout => \uart_tx_N_186_1\,
            ltout => \uart_tx_N_186_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNI2B741_0_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2219\,
            in3 => \N__2600\,
            lcout => \un1_M_count_q_ac0_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_1_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001111000"
        )
    port map (
            in0 => \N__2216\,
            in1 => \N__2733\,
            in2 => \N__2091\,
            in3 => \N__2748\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3192\,
            ce => 'H',
            sr => \N__2564\
        );

    \M_count_q_RNITRFR_3_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2189\,
            in2 => \_gnd_net_\,
            in3 => \N__2599\,
            lcout => OPEN,
            ltout => \un1_M_count_q_ac0_5_m2_0_a2_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_RNIF6FD2_1_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2666\,
            in1 => \N__2148\,
            in2 => \N__2114\,
            in3 => \N__2080\,
            lcout => \un1_M_count_q_ac0_5_m2_0_a2_3\,
            ltout => \un1_M_count_q_ac0_5_m2_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_4_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001101010"
        )
    port map (
            in0 => \N__2916\,
            in1 => \N__2734\,
            in2 => \N__2939\,
            in3 => \N__2749\,
            lcout => led_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3192\,
            ce => 'H',
            sr => \N__2564\
        );

    \click_dtct.M_last_q_RNIUTK51_0_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__2882\,
            in1 => \N__2858\,
            in2 => \N__2821\,
            in3 => \N__2779\,
            lcout => click_dtct_out8,
            ltout => \click_dtct_out8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_count_q_0_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011010101010"
        )
    port map (
            in0 => \N__2601\,
            in1 => \N__2732\,
            in2 => \N__2711\,
            in3 => \N__2667\,
            lcout => led_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3192\,
            ce => 'H',
            sr => \N__2564\
        );

    \btn_cond.M_ctr_q_0_LC_18_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2504\,
            in2 => \N__2519\,
            in3 => \N__2518\,
            lcout => \btn_cond.M_ctr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_27_0_\,
            carryout => \btn_cond.un1_M_ctr_q_cry_0\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_1_LC_18_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2486\,
            in2 => \_gnd_net_\,
            in3 => \N__2468\,
            lcout => \btn_cond.M_ctr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_0\,
            carryout => \btn_cond.un1_M_ctr_q_cry_1\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_2_LC_18_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2464\,
            in2 => \_gnd_net_\,
            in3 => \N__2444\,
            lcout => \btn_cond.M_ctr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_1\,
            carryout => \btn_cond.un1_M_ctr_q_cry_2\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_3_LC_18_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2436\,
            in2 => \_gnd_net_\,
            in3 => \N__2414\,
            lcout => \btn_cond.M_ctr_qZ0Z_3\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_2\,
            carryout => \btn_cond.un1_M_ctr_q_cry_3\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_4_LC_18_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2411\,
            in2 => \_gnd_net_\,
            in3 => \N__2393\,
            lcout => \btn_cond.M_ctr_qZ0Z_4\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_3\,
            carryout => \btn_cond.un1_M_ctr_q_cry_4\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_5_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3128\,
            in2 => \_gnd_net_\,
            in3 => \N__3110\,
            lcout => \btn_cond.M_ctr_qZ0Z_5\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_4\,
            carryout => \btn_cond.un1_M_ctr_q_cry_5\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_6_LC_18_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3107\,
            in2 => \_gnd_net_\,
            in3 => \N__3089\,
            lcout => \btn_cond.M_ctr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_5\,
            carryout => \btn_cond.un1_M_ctr_q_cry_6\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_7_LC_18_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3084\,
            in2 => \_gnd_net_\,
            in3 => \N__3059\,
            lcout => \btn_cond.M_ctr_qZ0Z_7\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_6\,
            carryout => \btn_cond.un1_M_ctr_q_cry_7\,
            clk => \N__3193\,
            ce => 'H',
            sr => \N__3143\
        );

    \btn_cond.M_ctr_q_8_LC_18_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3055\,
            in2 => \_gnd_net_\,
            in3 => \N__3035\,
            lcout => \btn_cond.M_ctr_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_28_0_\,
            carryout => \btn_cond.un1_M_ctr_q_cry_8\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_9_LC_18_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3032\,
            in2 => \_gnd_net_\,
            in3 => \N__3014\,
            lcout => \btn_cond.M_ctr_qZ0Z_9\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_8\,
            carryout => \btn_cond.un1_M_ctr_q_cry_9\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_10_LC_18_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3006\,
            in2 => \_gnd_net_\,
            in3 => \N__2984\,
            lcout => \btn_cond.M_ctr_qZ0Z_10\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_9\,
            carryout => \btn_cond.un1_M_ctr_q_cry_10\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_11_LC_18_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2981\,
            in2 => \_gnd_net_\,
            in3 => \N__2963\,
            lcout => \btn_cond.M_ctr_qZ0Z_11\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_10\,
            carryout => \btn_cond.un1_M_ctr_q_cry_11\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_12_LC_18_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2960\,
            in2 => \_gnd_net_\,
            in3 => \N__2942\,
            lcout => \btn_cond.M_ctr_qZ0Z_12\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_11\,
            carryout => \btn_cond.un1_M_ctr_q_cry_12\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_13_LC_18_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3355\,
            in2 => \_gnd_net_\,
            in3 => \N__3335\,
            lcout => \btn_cond.M_ctr_qZ0Z_13\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_12\,
            carryout => \btn_cond.un1_M_ctr_q_cry_13\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_14_LC_18_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3331\,
            in2 => \_gnd_net_\,
            in3 => \N__3308\,
            lcout => \btn_cond.M_ctr_qZ0Z_14\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_13\,
            carryout => \btn_cond.un1_M_ctr_q_cry_14\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_15_LC_18_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3304\,
            in2 => \_gnd_net_\,
            in3 => \N__3284\,
            lcout => \btn_cond.M_ctr_qZ0Z_15\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_14\,
            carryout => \btn_cond.un1_M_ctr_q_cry_15\,
            clk => \N__3194\,
            ce => 'H',
            sr => \N__3142\
        );

    \btn_cond.M_ctr_q_16_LC_18_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3276\,
            in2 => \_gnd_net_\,
            in3 => \N__3260\,
            lcout => \btn_cond.M_ctr_qZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_29_0_\,
            carryout => \btn_cond.un1_M_ctr_q_cry_16\,
            clk => \N__3196\,
            ce => 'H',
            sr => \N__3141\
        );

    \btn_cond.M_ctr_q_17_LC_18_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3255\,
            in2 => \_gnd_net_\,
            in3 => \N__3239\,
            lcout => \btn_cond.M_ctr_qZ0Z_17\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_16\,
            carryout => \btn_cond.un1_M_ctr_q_cry_17\,
            clk => \N__3196\,
            ce => 'H',
            sr => \N__3141\
        );

    \btn_cond.M_ctr_q_18_LC_18_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3236\,
            in2 => \_gnd_net_\,
            in3 => \N__3221\,
            lcout => \btn_cond.M_ctr_qZ0Z_18\,
            ltout => OPEN,
            carryin => \btn_cond.un1_M_ctr_q_cry_17\,
            carryout => \btn_cond.un1_M_ctr_q_cry_18\,
            clk => \N__3196\,
            ce => 'H',
            sr => \N__3141\
        );

    \btn_cond.M_ctr_q_19_LC_18_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3214\,
            in2 => \_gnd_net_\,
            in3 => \N__3218\,
            lcout => \btn_cond.M_ctr_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3196\,
            ce => 'H',
            sr => \N__3141\
        );
end \INTERFACE\;
